LIBRARY ieee;              
--USE ieee.std_logic_arith.all;                                 
USE ieee.std_logic_1164.all;  
USE ieee.numeric_std.all; 
USE ieee.std_logic_signed .all ;
USE ieee.std_logic_1164.std_ulogic;
------------------------------------------------------
ENTITY mining_hardware_var_tb IS
GENERIC	( 	  -- GENERIC funcion_hash

				  nonceL		   		: INTEGER	:= 32		;
				  
				  -- GENERIC generacion_nonce
				  
				  randL		   		: INTEGER	:= 12 		;
				  halfL  				: INTEGER	:= 6  	;  
				  sequL					: INTEGER	:= 20		;
				  twicL					: INTEGER	:= 24		;
				  
				  -- GENERIC comunicacion
				  
				  Convel    			: INTEGER  	:= 104	;  
			     Nvel      			: INTEGER  	:= 7		;
				  Conceros				: INTEGER  	:= 16		; 
				  Nceros					: INTEGER  	:= 5		;
				  Confinal				: INTEGER  	:= 208  	; 
				  Nfinal					: INTEGER  	:= 8		;
				  Conmitadvel 			: INTEGER  	:= 52  	;  
				  Nmitadvel      		: INTEGER  	:= 6		;
				  Conbits     			: INTEGER  	:= 7		;	  
				  Nbits					: INTEGER  	:= 3		;
				  Con512     			: INTEGER  	:= 511	;  
				  N512					: INTEGER  	:= 9		;
				  Conblock    			: INTEGER  	:= 16		;	  
				  Nblock					: INTEGER  	:= 5		;
				  Contransmision		: INTEGER  	:= 104  	;  
				  Ntransmision			: INTEGER  	:= 7		;
				  Conbits2    			: INTEGER  	:= 380	;  
				  Nbits2					: INTEGER  	:= 9		;
				  Xmax 					: INTEGER	:= 511	;
				  Ymax 					: INTEGER	:= 16		;
				  MAX_WIDTH			   : INTEGER	:= 380	;
				  Cont1     			: INTEGER	:= 100	;
				  Cont2		         : INTEGER 	:= 9		;
				  N1				      : INTEGER   := 10		;
				  N2			      	: INTEGER   := 4		;
				  Conad					: INTEGER	:= 100	;
				  Nad						: INTEGER	:= 10		);
END ENTITY;
------------------------------------------------------
ARCHITECTURE testbench_var_hw OF mining_hardware_var_tb IS 
SIGNAL  clk	               				:	STD_ULOGIC;
SIGNAL  rst, Rx, Tx							:	STD_ULOGIC;
--SIGNAL  entrada								:	STD_ULOGIC_VECTOR(1980 DOWNTO 0):="1100010110010000011001000000000100000000010000000001000000000101100111010011101101001100110101000011010100101101010101110101100111010011001101011001110100111011010000101101010101110100010011010000101101001101110100111011010101011101000110110100100011010001001101000010110101101011010011011101010101110100001011010010111101001000110101100111010110101101010101110100100011010000101101000100110101101011010010111101001000110101100111010001001101011010110100110111010010001101000010110100101111010001001101010101110100110111010010001101011010110100010011010111001101001010110100001011010010001101001100110100110111010111001101000100110100110011010110101101001010110100100011010011011101011010110101100111010100001101000100110100101011010010001101011010110100101111010010101101000010110100010011010010001101011010110100101011010110011101011100110100100011010011001101001101110101101011010111001101001100110100100011010111001101001101110101110011010001001101001101110100100011010000101101001101110101101011010111001101000100110100100011010101011101000100110101001111010110011101001000110100010011010000101101001000110100110111010111001101000010110100010011010010101101001000110100110111010010101101011001110100100011010001001101001101110101101011010000101101000100110101110011010000000011000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000101100000010000101111111111111111111111111111111111111111111";
--SIGNAL  entrada								:	STD_ULOGIC_VECTOR(1340 DOWNTO 0):="110000111001000001100100000000010000000001000000000100000000010100001101001000110101100011010001001101001000110101100011010001001101010100110101100011010001001101010100110100110011010001001101010100110100110011010111001101010100110100110011010111001101000010110100110011010111001101000010110101001011010111001101000010110101001011010010101101000010110101001011010010101101011010110101001011010010101101011010110100011011010010101101011010110100011011010101101101011010110100011011010101101101001110110100011011010101101101001110110101111011010101101101001110110101111011010000011101001110110101111011010000011101010001110100000000110000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000101000000010000001111111111111111111111111111111111111111111";
--SIGNAL  entrada								:	STD_ULOGIC_VECTOR(1340 DOWNTO 0):="110000011001000001100100000000010000000001000000000100000000010100001101001000110101100011010001001101001000110101100011010001001101010100110101100011010001001101010100110100110011010001001101010100110100110011010111001101010100110100110011010111001101000010110100110011010111001101000010110101001011010111001101000010110101001011010010101101000010110101001011010010101101011010110101001011010010101101011010110100011011010010101101011010110100011011010101101101011010110100011011010101101101001110110100011011010101101101001110110101111011010101101101001110110101111011010000011101001110110101111011010000011101010001110100000000110000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000101000000010000001111111111111111111111111111111111111111111";
SIGNAL  entrada								:	STD_ULOGIC_VECTOR(685 DOWNTO 0):="11000001100100000110010000000001000000000100000000010000000001010000110100100011010110001101000000001100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000111001111111111111111111111111";
--SIGNAL	i										: INTEGER :=1980;
--SIGNAL  i										:	INTEGER:=1340;
SIGNAL  i										:	INTEGER:=685;


BEGIN
	-------------- CLK GENERATION-------------------
	ClkGeneration: PROCESS
	BEGIN
		clk <= '0'; 
		WAIT FOR 10 ns;
		clk <= '1';
		WAIT FOR 10 ns;
	END PROCESS ClkGeneration;
	------------------------------------------------
	
	------- RESET GENERATION --------------------
	
	rstGeneration: PROCESS
	BEGIN		
		rst		<= '0' AFTER 10 ns,
						'1' AFTER 30 ns;
		WAIT FOR 100000 ms;
	END PROCESS rstGeneration;
	
	
	-------- Get hash signal in SHA block ------------
	
	serial: PROCESS
	BEGIN		
		
		FOR i IN 685 DOWNTO 0 LOOP
		Rx		<= entrada(i);		
		WAIT FOR 2.14 us;
		END LOOP;
	END PROCESS serial;
	
	
	-- Component Instantiation DUT (Device Under Test)
	
	ModuleDUT_hw: ENTITY work.mining_hardware_var
	GENERIC	MAP( 	nonceL		   	=>	nonceL,
						
						randL					=> randL,	 
						halfL  	  			=> halfL,
						sequL					=> sequL,
						twicL					=> twicL,
						
						Convel    		   => Convel,  
					   Nvel      			=> Nvel,
					   Conceros				=> Conceros, 
					   Nceros				=> Nceros,
					   Confinal				=> Confinal, 
					   Nfinal				=> Nfinal,
					   Conmitadvel 		=> Conmitadvel, 
					   Nmitadvel      	=> Nmitadvel,
					   Conbits     		=> Conbits,  
					   Nbits					=> Nbits,
					   Con512     			=> Con512,  
					   N512					=> N512,
					   Conblock    		=> Conblock,  
					   Nblock				=> Nblock,
					   Contransmision		=> Contransmision, 
					   Ntransmision		=> Ntransmision,
					   Conbits2    		=> Conbits2,  
					   Nbits2				=> Nbits2,
					   Xmax 					=> Xmax,
					   Ymax 					=> Ymax,
					   MAX_WIDTH			=> MAX_WIDTH,
						Cont1 				=> Cont1,
						Cont2					=> Cont2,
						N1						=> N1,
						N2						=> N2,
						Conad					=> Conad,
						Nad					=> Nad
					)
	PORT	  MAP ( clk	    	=>		clk,
					  rst			=>		rst,
					  Rx        =>    Rx,
					  Tx			=> 	Tx
					 );
					 
	--------------------------------------------------					  
END ARCHITECTURE testbench_var_hw;	