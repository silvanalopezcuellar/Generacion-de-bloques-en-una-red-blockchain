LIBRARY IEEE;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
----------------------------------
ENTITY Output_sel IS
	GENERIC  ( BitsNonce				:	INTEGER := 32);   
	PORT		( clk						:	IN		STD_ULOGIC;
				  rst						:	IN 	STD_ULOGIC;
				  ceros_ok				:	IN		STD_ULOGIC_VECTOR(15 DOWNTO 0);
				  enable					:	IN		STD_ULOGIC;
				  output0				:	IN		STD_ULOGIC_VECTOR(255 DOWNTO 0);
				  output1				:	IN		STD_ULOGIC_VECTOR(255 DOWNTO 0);
				  output2				:	IN		STD_ULOGIC_VECTOR(255 DOWNTO 0);
				  output3				:	IN		STD_ULOGIC_VECTOR(255 DOWNTO 0);
				  output4				:	IN		STD_ULOGIC_VECTOR(255 DOWNTO 0);
				  output5				:	IN		STD_ULOGIC_VECTOR(255 DOWNTO 0);
				  output6				:	IN		STD_ULOGIC_VECTOR(255 DOWNTO 0);
				  output7				:	IN		STD_ULOGIC_VECTOR(255 DOWNTO 0);
				  output8				:	IN		STD_ULOGIC_VECTOR(255 DOWNTO 0);
				  output9				:	IN		STD_ULOGIC_VECTOR(255 DOWNTO 0);
				  outputA				:	IN		STD_ULOGIC_VECTOR(255 DOWNTO 0);
				  outputB				:	IN		STD_ULOGIC_VECTOR(255 DOWNTO 0);
				  outputC				:	IN		STD_ULOGIC_VECTOR(255 DOWNTO 0);
				  outputD				:	IN		STD_ULOGIC_VECTOR(255 DOWNTO 0);
				  outputE				:	IN		STD_ULOGIC_VECTOR(255 DOWNTO 0);
				  outputF				:	IN		STD_ULOGIC_VECTOR(255 DOWNTO 0);
				  nonce0					:	IN		STD_ULOGIC_VECTOR(BitsNonce-1 DOWNTO 0);
				  nonce1					:	IN		STD_ULOGIC_VECTOR(BitsNonce-1 DOWNTO 0);
				  nonce2					:	IN		STD_ULOGIC_VECTOR(BitsNonce-1 DOWNTO 0);
				  nonce3					:	IN		STD_ULOGIC_VECTOR(BitsNonce-1 DOWNTO 0);
				  nonce4					:	IN		STD_ULOGIC_VECTOR(BitsNonce-1 DOWNTO 0);
				  nonce5					:	IN		STD_ULOGIC_VECTOR(BitsNonce-1 DOWNTO 0);
				  nonce6					:	IN		STD_ULOGIC_VECTOR(BitsNonce-1 DOWNTO 0);
				  nonce7					:	IN		STD_ULOGIC_VECTOR(BitsNonce-1 DOWNTO 0);
				  nonce8					:	IN		STD_ULOGIC_VECTOR(BitsNonce-1 DOWNTO 0);
				  nonce9					:	IN		STD_ULOGIC_VECTOR(BitsNonce-1 DOWNTO 0);
				  nonceA					:	IN		STD_ULOGIC_VECTOR(BitsNonce-1 DOWNTO 0);
				  nonceB					:	IN		STD_ULOGIC_VECTOR(BitsNonce-1 DOWNTO 0);
				  nonceC					:	IN		STD_ULOGIC_VECTOR(BitsNonce-1 DOWNTO 0);
				  nonceD					:	IN		STD_ULOGIC_VECTOR(BitsNonce-1 DOWNTO 0);
				  nonceE					:	IN		STD_ULOGIC_VECTOR(BitsNonce-1 DOWNTO 0);
				  nonceF					:	IN		STD_ULOGIC_VECTOR(BitsNonce-1 DOWNTO 0);
				  salida_final			:	OUT   STD_ULOGIC_VECTOR(287 DOWNTO 0));
END ENTITY;
---------------------------------- 

----------------------------------
ARCHITECTURE Output_selArchh OF Output_sel IS
	SIGNAL	registro_final		:	STD_ULOGIC_VECTOR(287 DOWNTO 0); 
BEGIN
			SALida_final <= registro_final;
	PROCESS(clk,rst, enable)
	BEGIN
		IF(rst = '0') THEN
			registro_final <= (OTHERS => '0');
		ELSIF(RISING_EDGE(clk)) THEN
			IF( (enable = '1' ) ) THEN
			registro_final(0) <= (nonce0(0) AND ceros_ok(0)) OR (nonce1(0) AND ceros_ok(1)) OR (nonce2(0) AND ceros_ok(2)) OR (nonce3(0) AND ceros_ok(3)) OR (nonce4(0) AND ceros_ok(4)) OR (nonce5(0) AND ceros_ok(5)) OR (nonce6(0) AND ceros_ok(6)) OR (nonce7(0) AND ceros_ok(7))OR (nonce8(0) AND ceros_ok(8))OR (nonce9(0) AND ceros_ok(9)) OR (nonceA(0) AND ceros_ok(10)) OR (nonceB(0) AND ceros_ok(11)) OR (nonceC(0) AND ceros_ok(12)) OR (nonceD(0) AND ceros_ok(13)) OR (nonceE(0) AND ceros_ok(14)) OR (nonceF(0) AND ceros_ok(15));
			registro_final(1) <= (nonce0(1) AND ceros_ok(0)) OR (nonce1(1) AND ceros_ok(1)) OR (nonce2(1) AND ceros_ok(2)) OR (nonce3(1) AND ceros_ok(3)) OR (nonce4(1) AND ceros_ok(4)) OR (nonce5(1) AND ceros_ok(5)) OR (nonce6(1) AND ceros_ok(6)) OR (nonce7(1) AND ceros_ok(7))OR (nonce8(1) AND ceros_ok(8))OR (nonce9(1) AND ceros_ok(9)) OR (nonceA(1) AND ceros_ok(10)) OR (nonceB(1) AND ceros_ok(11)) OR (nonceC(1) AND ceros_ok(12)) OR (nonceD(1) AND ceros_ok(13)) OR (nonceE(1) AND ceros_ok(14)) OR (nonceF(1) AND ceros_ok(15));
			registro_final(2) <= (nonce0(2) AND ceros_ok(0)) OR (nonce1(2) AND ceros_ok(1)) OR (nonce2(2) AND ceros_ok(2)) OR (nonce3(2) AND ceros_ok(3)) OR (nonce4(2) AND ceros_ok(4)) OR (nonce5(2) AND ceros_ok(5)) OR (nonce6(2) AND ceros_ok(6)) OR (nonce7(2) AND ceros_ok(7))OR (nonce8(2) AND ceros_ok(8))OR (nonce9(2) AND ceros_ok(9)) OR (nonceA(2) AND ceros_ok(10)) OR (nonceB(2) AND ceros_ok(11)) OR (nonceC(2) AND ceros_ok(12)) OR (nonceD(2) AND ceros_ok(13)) OR (nonceE(2) AND ceros_ok(14)) OR (nonceF(2) AND ceros_ok(15));
			registro_final(3) <= (nonce0(3) AND ceros_ok(0)) OR (nonce1(3) AND ceros_ok(1)) OR (nonce2(3) AND ceros_ok(2)) OR (nonce3(3) AND ceros_ok(3)) OR (nonce4(3) AND ceros_ok(4)) OR (nonce5(3) AND ceros_ok(5)) OR (nonce6(3) AND ceros_ok(6)) OR (nonce7(3) AND ceros_ok(7))OR (nonce8(3) AND ceros_ok(8))OR (nonce9(3) AND ceros_ok(9)) OR (nonceA(3) AND ceros_ok(10)) OR (nonceB(3) AND ceros_ok(11)) OR (nonceC(3) AND ceros_ok(12)) OR (nonceD(3) AND ceros_ok(13)) OR (nonceE(3) AND ceros_ok(14)) OR (nonceF(3) AND ceros_ok(15));
			registro_final(4) <= (nonce0(4) AND ceros_ok(0)) OR (nonce1(4) AND ceros_ok(1)) OR (nonce2(4) AND ceros_ok(2)) OR (nonce3(4) AND ceros_ok(3)) OR (nonce4(4) AND ceros_ok(4)) OR (nonce5(4) AND ceros_ok(5)) OR (nonce6(4) AND ceros_ok(6)) OR (nonce7(4) AND ceros_ok(7))OR (nonce8(4) AND ceros_ok(8))OR (nonce9(4) AND ceros_ok(9)) OR (nonceA(4) AND ceros_ok(10)) OR (nonceB(4) AND ceros_ok(11)) OR (nonceC(4) AND ceros_ok(12)) OR (nonceD(4) AND ceros_ok(13)) OR (nonceE(4) AND ceros_ok(14)) OR (nonceF(4) AND ceros_ok(15));
			registro_final(5) <= (nonce0(5) AND ceros_ok(0)) OR (nonce1(5) AND ceros_ok(1)) OR (nonce2(5) AND ceros_ok(2)) OR (nonce3(5) AND ceros_ok(3)) OR (nonce4(5) AND ceros_ok(4)) OR (nonce5(5) AND ceros_ok(5)) OR (nonce6(5) AND ceros_ok(6)) OR (nonce7(5) AND ceros_ok(7))OR (nonce8(5) AND ceros_ok(8))OR (nonce9(5) AND ceros_ok(9)) OR (nonceA(5) AND ceros_ok(10)) OR (nonceB(5) AND ceros_ok(11)) OR (nonceC(5) AND ceros_ok(12)) OR (nonceD(5) AND ceros_ok(13)) OR (nonceE(5) AND ceros_ok(14)) OR (nonceF(5) AND ceros_ok(15));
			registro_final(6) <= (nonce0(6) AND ceros_ok(0)) OR (nonce1(6) AND ceros_ok(1)) OR (nonce2(6) AND ceros_ok(2)) OR (nonce3(6) AND ceros_ok(3)) OR (nonce4(6) AND ceros_ok(4)) OR (nonce5(6) AND ceros_ok(5)) OR (nonce6(6) AND ceros_ok(6)) OR (nonce7(6) AND ceros_ok(7))OR (nonce8(6) AND ceros_ok(8))OR (nonce9(6) AND ceros_ok(9)) OR (nonceA(6) AND ceros_ok(10)) OR (nonceB(6) AND ceros_ok(11)) OR (nonceC(6) AND ceros_ok(12)) OR (nonceD(6) AND ceros_ok(13)) OR (nonceE(6) AND ceros_ok(14)) OR (nonceF(6) AND ceros_ok(15));
			registro_final(7) <= (nonce0(7) AND ceros_ok(0)) OR (nonce1(7) AND ceros_ok(1)) OR (nonce2(7) AND ceros_ok(2)) OR (nonce3(7) AND ceros_ok(3)) OR (nonce4(7) AND ceros_ok(4)) OR (nonce5(7) AND ceros_ok(5)) OR (nonce6(7) AND ceros_ok(6)) OR (nonce7(7) AND ceros_ok(7))OR (nonce8(7) AND ceros_ok(8))OR (nonce9(7) AND ceros_ok(9)) OR (nonceA(7) AND ceros_ok(10)) OR (nonceB(7) AND ceros_ok(11)) OR (nonceC(7) AND ceros_ok(12)) OR (nonceD(7) AND ceros_ok(13)) OR (nonceE(7) AND ceros_ok(14)) OR (nonceF(7) AND ceros_ok(15));
			registro_final(8) <= (nonce0(8) AND ceros_ok(0)) OR (nonce1(8) AND ceros_ok(1)) OR (nonce2(8) AND ceros_ok(2)) OR (nonce3(8) AND ceros_ok(3)) OR (nonce4(8) AND ceros_ok(4)) OR (nonce5(8) AND ceros_ok(5)) OR (nonce6(8) AND ceros_ok(6)) OR (nonce7(8) AND ceros_ok(7))OR (nonce8(8) AND ceros_ok(8))OR (nonce9(8) AND ceros_ok(9)) OR (nonceA(8) AND ceros_ok(10)) OR (nonceB(8) AND ceros_ok(11)) OR (nonceC(8) AND ceros_ok(12)) OR (nonceD(8) AND ceros_ok(13)) OR (nonceE(8) AND ceros_ok(14)) OR (nonceF(8) AND ceros_ok(15));
			registro_final(9) <= (nonce0(9) AND ceros_ok(0)) OR (nonce1(9) AND ceros_ok(1)) OR (nonce2(9) AND ceros_ok(2)) OR (nonce3(9) AND ceros_ok(3)) OR (nonce4(9) AND ceros_ok(4)) OR (nonce5(9) AND ceros_ok(5)) OR (nonce6(9) AND ceros_ok(6)) OR (nonce7(9) AND ceros_ok(7))OR (nonce8(9) AND ceros_ok(8))OR (nonce9(9) AND ceros_ok(9)) OR (nonceA(9) AND ceros_ok(10)) OR (nonceB(9) AND ceros_ok(11)) OR (nonceC(9) AND ceros_ok(12)) OR (nonceD(9) AND ceros_ok(13)) OR (nonceE(9) AND ceros_ok(14)) OR (nonceF(9) AND ceros_ok(15));
			registro_final(10) <= (nonce0(10) AND ceros_ok(0)) OR (nonce1(10) AND ceros_ok(1)) OR (nonce2(10) AND ceros_ok(2)) OR (nonce3(10) AND ceros_ok(3)) OR (nonce4(10) AND ceros_ok(4)) OR (nonce5(10) AND ceros_ok(5)) OR (nonce6(10) AND ceros_ok(6)) OR (nonce7(10) AND ceros_ok(7))OR (nonce8(10) AND ceros_ok(8))OR (nonce9(10) AND ceros_ok(9)) OR (nonceA(10) AND ceros_ok(10)) OR (nonceB(10) AND ceros_ok(11)) OR (nonceC(10) AND ceros_ok(12)) OR (nonceD(10) AND ceros_ok(13)) OR (nonceE(10) AND ceros_ok(14)) OR (nonceF(10) AND ceros_ok(15));
			registro_final(11) <= (nonce0(11) AND ceros_ok(0)) OR (nonce1(11) AND ceros_ok(1)) OR (nonce2(11) AND ceros_ok(2)) OR (nonce3(11) AND ceros_ok(3)) OR (nonce4(11) AND ceros_ok(4)) OR (nonce5(11) AND ceros_ok(5)) OR (nonce6(11) AND ceros_ok(6)) OR (nonce7(11) AND ceros_ok(7))OR (nonce8(11) AND ceros_ok(8))OR (nonce9(11) AND ceros_ok(9)) OR (nonceA(11) AND ceros_ok(10)) OR (nonceB(11) AND ceros_ok(11)) OR (nonceC(11) AND ceros_ok(12)) OR (nonceD(11) AND ceros_ok(13)) OR (nonceE(11) AND ceros_ok(14)) OR (nonceF(11) AND ceros_ok(15));
			registro_final(12) <= (nonce0(12) AND ceros_ok(0)) OR (nonce1(12) AND ceros_ok(1)) OR (nonce2(12) AND ceros_ok(2)) OR (nonce3(12) AND ceros_ok(3)) OR (nonce4(12) AND ceros_ok(4)) OR (nonce5(12) AND ceros_ok(5)) OR (nonce6(12) AND ceros_ok(6)) OR (nonce7(12) AND ceros_ok(7))OR (nonce8(12) AND ceros_ok(8))OR (nonce9(12) AND ceros_ok(9)) OR (nonceA(12) AND ceros_ok(10)) OR (nonceB(12) AND ceros_ok(11)) OR (nonceC(12) AND ceros_ok(12)) OR (nonceD(12) AND ceros_ok(13)) OR (nonceE(12) AND ceros_ok(14)) OR (nonceF(12) AND ceros_ok(15));
			registro_final(13) <= (nonce0(13) AND ceros_ok(0)) OR (nonce1(13) AND ceros_ok(1)) OR (nonce2(13) AND ceros_ok(2)) OR (nonce3(13) AND ceros_ok(3)) OR (nonce4(13) AND ceros_ok(4)) OR (nonce5(13) AND ceros_ok(5)) OR (nonce6(13) AND ceros_ok(6)) OR (nonce7(13) AND ceros_ok(7))OR (nonce8(13) AND ceros_ok(8))OR (nonce9(13) AND ceros_ok(9)) OR (nonceA(13) AND ceros_ok(10)) OR (nonceB(13) AND ceros_ok(11)) OR (nonceC(13) AND ceros_ok(12)) OR (nonceD(13) AND ceros_ok(13)) OR (nonceE(13) AND ceros_ok(14)) OR (nonceF(13) AND ceros_ok(15));
			registro_final(14) <= (nonce0(14) AND ceros_ok(0)) OR (nonce1(14) AND ceros_ok(1)) OR (nonce2(14) AND ceros_ok(2)) OR (nonce3(14) AND ceros_ok(3)) OR (nonce4(14) AND ceros_ok(4)) OR (nonce5(14) AND ceros_ok(5)) OR (nonce6(14) AND ceros_ok(6)) OR (nonce7(14) AND ceros_ok(7))OR (nonce8(14) AND ceros_ok(8))OR (nonce9(14) AND ceros_ok(9)) OR (nonceA(14) AND ceros_ok(10)) OR (nonceB(14) AND ceros_ok(11)) OR (nonceC(14) AND ceros_ok(12)) OR (nonceD(14) AND ceros_ok(13)) OR (nonceE(14) AND ceros_ok(14)) OR (nonceF(14) AND ceros_ok(15));
			registro_final(15) <= (nonce0(15) AND ceros_ok(0)) OR (nonce1(15) AND ceros_ok(1)) OR (nonce2(15) AND ceros_ok(2)) OR (nonce3(15) AND ceros_ok(3)) OR (nonce4(15) AND ceros_ok(4)) OR (nonce5(15) AND ceros_ok(5)) OR (nonce6(15) AND ceros_ok(6)) OR (nonce7(15) AND ceros_ok(7))OR (nonce8(15) AND ceros_ok(8))OR (nonce9(15) AND ceros_ok(9)) OR (nonceA(15) AND ceros_ok(10)) OR (nonceB(15) AND ceros_ok(11)) OR (nonceC(15) AND ceros_ok(12)) OR (nonceD(15) AND ceros_ok(13)) OR (nonceE(15) AND ceros_ok(14)) OR (nonceF(15) AND ceros_ok(15));
			registro_final(16) <= (nonce0(16) AND ceros_ok(0)) OR (nonce1(16) AND ceros_ok(1)) OR (nonce2(16) AND ceros_ok(2)) OR (nonce3(16) AND ceros_ok(3)) OR (nonce4(16) AND ceros_ok(4)) OR (nonce5(16) AND ceros_ok(5)) OR (nonce6(16) AND ceros_ok(6)) OR (nonce7(16) AND ceros_ok(7))OR (nonce8(16) AND ceros_ok(8))OR (nonce9(16) AND ceros_ok(9)) OR (nonceA(16) AND ceros_ok(10)) OR (nonceB(16) AND ceros_ok(11)) OR (nonceC(16) AND ceros_ok(12)) OR (nonceD(16) AND ceros_ok(13)) OR (nonceE(16) AND ceros_ok(14)) OR (nonceF(16) AND ceros_ok(15));
			registro_final(17) <= (nonce0(17) AND ceros_ok(0)) OR (nonce1(17) AND ceros_ok(1)) OR (nonce2(17) AND ceros_ok(2)) OR (nonce3(17) AND ceros_ok(3)) OR (nonce4(17) AND ceros_ok(4)) OR (nonce5(17) AND ceros_ok(5)) OR (nonce6(17) AND ceros_ok(6)) OR (nonce7(17) AND ceros_ok(7))OR (nonce8(17) AND ceros_ok(8))OR (nonce9(17) AND ceros_ok(9)) OR (nonceA(17) AND ceros_ok(10)) OR (nonceB(17) AND ceros_ok(11)) OR (nonceC(17) AND ceros_ok(12)) OR (nonceD(17) AND ceros_ok(13)) OR (nonceE(17) AND ceros_ok(14)) OR (nonceF(17) AND ceros_ok(15));
			registro_final(18) <= (nonce0(18) AND ceros_ok(0)) OR (nonce1(18) AND ceros_ok(1)) OR (nonce2(18) AND ceros_ok(2)) OR (nonce3(18) AND ceros_ok(3)) OR (nonce4(18) AND ceros_ok(4)) OR (nonce5(18) AND ceros_ok(5)) OR (nonce6(18) AND ceros_ok(6)) OR (nonce7(18) AND ceros_ok(7))OR (nonce8(18) AND ceros_ok(8))OR (nonce9(18) AND ceros_ok(9)) OR (nonceA(18) AND ceros_ok(10)) OR (nonceB(18) AND ceros_ok(11)) OR (nonceC(18) AND ceros_ok(12)) OR (nonceD(18) AND ceros_ok(13)) OR (nonceE(18) AND ceros_ok(14)) OR (nonceF(18) AND ceros_ok(15));
			registro_final(19) <= (nonce0(19) AND ceros_ok(0)) OR (nonce1(19) AND ceros_ok(1)) OR (nonce2(19) AND ceros_ok(2)) OR (nonce3(19) AND ceros_ok(3)) OR (nonce4(19) AND ceros_ok(4)) OR (nonce5(19) AND ceros_ok(5)) OR (nonce6(19) AND ceros_ok(6)) OR (nonce7(19) AND ceros_ok(7))OR (nonce8(19) AND ceros_ok(8))OR (nonce9(19) AND ceros_ok(9)) OR (nonceA(19) AND ceros_ok(10)) OR (nonceB(19) AND ceros_ok(11)) OR (nonceC(19) AND ceros_ok(12)) OR (nonceD(19) AND ceros_ok(13)) OR (nonceE(19) AND ceros_ok(14)) OR (nonceF(19) AND ceros_ok(15));
			registro_final(20) <= (nonce0(20) AND ceros_ok(0)) OR (nonce1(20) AND ceros_ok(1)) OR (nonce2(20) AND ceros_ok(2)) OR (nonce3(20) AND ceros_ok(3)) OR (nonce4(20) AND ceros_ok(4)) OR (nonce5(20) AND ceros_ok(5)) OR (nonce6(20) AND ceros_ok(6)) OR (nonce7(20) AND ceros_ok(7))OR (nonce8(20) AND ceros_ok(8))OR (nonce9(20) AND ceros_ok(9)) OR (nonceA(20) AND ceros_ok(10)) OR (nonceB(20) AND ceros_ok(11)) OR (nonceC(20) AND ceros_ok(12)) OR (nonceD(20) AND ceros_ok(13)) OR (nonceE(20) AND ceros_ok(14)) OR (nonceF(20) AND ceros_ok(15));
			registro_final(21) <= (nonce0(21) AND ceros_ok(0)) OR (nonce1(21) AND ceros_ok(1)) OR (nonce2(21) AND ceros_ok(2)) OR (nonce3(21) AND ceros_ok(3)) OR (nonce4(21) AND ceros_ok(4)) OR (nonce5(21) AND ceros_ok(5)) OR (nonce6(21) AND ceros_ok(6)) OR (nonce7(21) AND ceros_ok(7))OR (nonce8(21) AND ceros_ok(8))OR (nonce9(21) AND ceros_ok(9)) OR (nonceA(21) AND ceros_ok(10)) OR (nonceB(21) AND ceros_ok(11)) OR (nonceC(21) AND ceros_ok(12)) OR (nonceD(21) AND ceros_ok(13)) OR (nonceE(21) AND ceros_ok(14)) OR (nonceF(21) AND ceros_ok(15));
			registro_final(22) <= (nonce0(22) AND ceros_ok(0)) OR (nonce1(22) AND ceros_ok(1)) OR (nonce2(22) AND ceros_ok(2)) OR (nonce3(22) AND ceros_ok(3)) OR (nonce4(22) AND ceros_ok(4)) OR (nonce5(22) AND ceros_ok(5)) OR (nonce6(22) AND ceros_ok(6)) OR (nonce7(22) AND ceros_ok(7))OR (nonce8(22) AND ceros_ok(8))OR (nonce9(22) AND ceros_ok(9)) OR (nonceA(22) AND ceros_ok(10)) OR (nonceB(22) AND ceros_ok(11)) OR (nonceC(22) AND ceros_ok(12)) OR (nonceD(22) AND ceros_ok(13)) OR (nonceE(22) AND ceros_ok(14)) OR (nonceF(22) AND ceros_ok(15));
			registro_final(23) <= (nonce0(23) AND ceros_ok(0)) OR (nonce1(23) AND ceros_ok(1)) OR (nonce2(23) AND ceros_ok(2)) OR (nonce3(23) AND ceros_ok(3)) OR (nonce4(23) AND ceros_ok(4)) OR (nonce5(23) AND ceros_ok(5)) OR (nonce6(23) AND ceros_ok(6)) OR (nonce7(23) AND ceros_ok(7))OR (nonce8(23) AND ceros_ok(8))OR (nonce9(23) AND ceros_ok(9)) OR (nonceA(23) AND ceros_ok(10)) OR (nonceB(23) AND ceros_ok(11)) OR (nonceC(23) AND ceros_ok(12)) OR (nonceD(23) AND ceros_ok(13)) OR (nonceE(23) AND ceros_ok(14)) OR (nonceF(23) AND ceros_ok(15));
			registro_final(24) <= (nonce0(24) AND ceros_ok(0)) OR (nonce1(24) AND ceros_ok(1)) OR (nonce2(24) AND ceros_ok(2)) OR (nonce3(24) AND ceros_ok(3)) OR (nonce4(24) AND ceros_ok(4)) OR (nonce5(24) AND ceros_ok(5)) OR (nonce6(24) AND ceros_ok(6)) OR (nonce7(24) AND ceros_ok(7))OR (nonce8(24) AND ceros_ok(8))OR (nonce9(24) AND ceros_ok(9)) OR (nonceA(24) AND ceros_ok(10)) OR (nonceB(24) AND ceros_ok(11)) OR (nonceC(24) AND ceros_ok(12)) OR (nonceD(24) AND ceros_ok(13)) OR (nonceE(24) AND ceros_ok(14)) OR (nonceF(24) AND ceros_ok(15));
			registro_final(25) <= (nonce0(25) AND ceros_ok(0)) OR (nonce1(25) AND ceros_ok(1)) OR (nonce2(25) AND ceros_ok(2)) OR (nonce3(25) AND ceros_ok(3)) OR (nonce4(25) AND ceros_ok(4)) OR (nonce5(25) AND ceros_ok(5)) OR (nonce6(25) AND ceros_ok(6)) OR (nonce7(25) AND ceros_ok(7))OR (nonce8(25) AND ceros_ok(8))OR (nonce9(25) AND ceros_ok(9)) OR (nonceA(25) AND ceros_ok(10)) OR (nonceB(25) AND ceros_ok(11)) OR (nonceC(25) AND ceros_ok(12)) OR (nonceD(25) AND ceros_ok(13)) OR (nonceE(25) AND ceros_ok(14)) OR (nonceF(25) AND ceros_ok(15));
			registro_final(26) <= (nonce0(26) AND ceros_ok(0)) OR (nonce1(26) AND ceros_ok(1)) OR (nonce2(26) AND ceros_ok(2)) OR (nonce3(26) AND ceros_ok(3)) OR (nonce4(26) AND ceros_ok(4)) OR (nonce5(26) AND ceros_ok(5)) OR (nonce6(26) AND ceros_ok(6)) OR (nonce7(26) AND ceros_ok(7))OR (nonce8(26) AND ceros_ok(8))OR (nonce9(26) AND ceros_ok(9)) OR (nonceA(26) AND ceros_ok(10)) OR (nonceB(26) AND ceros_ok(11)) OR (nonceC(26) AND ceros_ok(12)) OR (nonceD(26) AND ceros_ok(13)) OR (nonceE(26) AND ceros_ok(14)) OR (nonceF(26) AND ceros_ok(15));
			registro_final(27) <= (nonce0(27) AND ceros_ok(0)) OR (nonce1(27) AND ceros_ok(1)) OR (nonce2(27) AND ceros_ok(2)) OR (nonce3(27) AND ceros_ok(3)) OR (nonce4(27) AND ceros_ok(4)) OR (nonce5(27) AND ceros_ok(5)) OR (nonce6(27) AND ceros_ok(6)) OR (nonce7(27) AND ceros_ok(7))OR (nonce8(27) AND ceros_ok(8))OR (nonce9(27) AND ceros_ok(9)) OR (nonceA(27) AND ceros_ok(10)) OR (nonceB(27) AND ceros_ok(11)) OR (nonceC(27) AND ceros_ok(12)) OR (nonceD(27) AND ceros_ok(13)) OR (nonceE(27) AND ceros_ok(14)) OR (nonceF(27) AND ceros_ok(15));
			registro_final(28) <= (nonce0(28) AND ceros_ok(0)) OR (nonce1(28) AND ceros_ok(1)) OR (nonce2(28) AND ceros_ok(2)) OR (nonce3(28) AND ceros_ok(3)) OR (nonce4(28) AND ceros_ok(4)) OR (nonce5(28) AND ceros_ok(5)) OR (nonce6(28) AND ceros_ok(6)) OR (nonce7(28) AND ceros_ok(7))OR (nonce8(28) AND ceros_ok(8))OR (nonce9(28) AND ceros_ok(9)) OR (nonceA(28) AND ceros_ok(10)) OR (nonceB(28) AND ceros_ok(11)) OR (nonceC(28) AND ceros_ok(12)) OR (nonceD(28) AND ceros_ok(13)) OR (nonceE(28) AND ceros_ok(14)) OR (nonceF(28) AND ceros_ok(15));
			registro_final(29) <= (nonce0(29) AND ceros_ok(0)) OR (nonce1(29) AND ceros_ok(1)) OR (nonce2(29) AND ceros_ok(2)) OR (nonce3(29) AND ceros_ok(3)) OR (nonce4(29) AND ceros_ok(4)) OR (nonce5(29) AND ceros_ok(5)) OR (nonce6(29) AND ceros_ok(6)) OR (nonce7(29) AND ceros_ok(7))OR (nonce8(29) AND ceros_ok(8))OR (nonce9(29) AND ceros_ok(9)) OR (nonceA(29) AND ceros_ok(10)) OR (nonceB(29) AND ceros_ok(11)) OR (nonceC(29) AND ceros_ok(12)) OR (nonceD(29) AND ceros_ok(13)) OR (nonceE(29) AND ceros_ok(14)) OR (nonceF(29) AND ceros_ok(15));
			registro_final(30) <= (nonce0(30) AND ceros_ok(0)) OR (nonce1(30) AND ceros_ok(1)) OR (nonce2(30) AND ceros_ok(2)) OR (nonce3(30) AND ceros_ok(3)) OR (nonce4(30) AND ceros_ok(4)) OR (nonce5(30) AND ceros_ok(5)) OR (nonce6(30) AND ceros_ok(6)) OR (nonce7(30) AND ceros_ok(7))OR (nonce8(30) AND ceros_ok(8))OR (nonce9(30) AND ceros_ok(9)) OR (nonceA(30) AND ceros_ok(10)) OR (nonceB(30) AND ceros_ok(11)) OR (nonceC(30) AND ceros_ok(12)) OR (nonceD(30) AND ceros_ok(13)) OR (nonceE(30) AND ceros_ok(14)) OR (nonceF(30) AND ceros_ok(15));
			registro_final(31) <= (nonce0(31) AND ceros_ok(0)) OR (nonce1(31) AND ceros_ok(1)) OR (nonce2(31) AND ceros_ok(2)) OR (nonce3(31) AND ceros_ok(3)) OR (nonce4(31) AND ceros_ok(4)) OR (nonce5(31) AND ceros_ok(5)) OR (nonce6(31) AND ceros_ok(6)) OR (nonce7(31) AND ceros_ok(7))OR (nonce8(31) AND ceros_ok(8))OR (nonce9(31) AND ceros_ok(9)) OR (nonceA(31) AND ceros_ok(10)) OR (nonceB(31) AND ceros_ok(11)) OR (nonceC(31) AND ceros_ok(12)) OR (nonceD(31) AND ceros_ok(13)) OR (nonceE(31) AND ceros_ok(14)) OR (nonceF(31) AND ceros_ok(15));
			registro_final(32) <= (output0(0) AND ceros_ok(0)) OR (output1(0) AND ceros_ok(1)) OR (output2(0) AND ceros_ok(2)) OR (output3(0) AND ceros_ok(3)) OR (output4(0) AND ceros_ok(4)) OR (output5(0) AND ceros_ok(5)) OR (output6(0) AND ceros_ok(6)) OR (output7(0) AND ceros_ok(7))OR (output8(0) AND ceros_ok(8))OR (output9(0) AND ceros_ok(9)) OR (outputA(0) AND ceros_ok(10)) OR (outputB(0) AND ceros_ok(11)) OR (outputC(0) AND ceros_ok(12)) OR (outputD(0) AND ceros_ok(13)) OR (outputE(0) AND ceros_ok(14)) OR (outputF(0) AND ceros_ok(15));
			registro_final(33) <= (output0(1) AND ceros_ok(0)) OR (output1(1) AND ceros_ok(1)) OR (output2(1) AND ceros_ok(2)) OR (output3(1) AND ceros_ok(3)) OR (output4(1) AND ceros_ok(4)) OR (output5(1) AND ceros_ok(5)) OR (output6(1) AND ceros_ok(6)) OR (output7(1) AND ceros_ok(7))OR (output8(1) AND ceros_ok(8))OR (output9(1) AND ceros_ok(9)) OR (outputA(1) AND ceros_ok(10)) OR (outputB(1) AND ceros_ok(11)) OR (outputC(1) AND ceros_ok(12)) OR (outputD(1) AND ceros_ok(13)) OR (outputE(1) AND ceros_ok(14)) OR (outputF(1) AND ceros_ok(15));
			registro_final(34) <= (output0(2) AND ceros_ok(0)) OR (output1(2) AND ceros_ok(1)) OR (output2(2) AND ceros_ok(2)) OR (output3(2) AND ceros_ok(3)) OR (output4(2) AND ceros_ok(4)) OR (output5(2) AND ceros_ok(5)) OR (output6(2) AND ceros_ok(6)) OR (output7(2) AND ceros_ok(7))OR (output8(2) AND ceros_ok(8))OR (output9(2) AND ceros_ok(9)) OR (outputA(2) AND ceros_ok(10)) OR (outputB(2) AND ceros_ok(11)) OR (outputC(2) AND ceros_ok(12)) OR (outputD(2) AND ceros_ok(13)) OR (outputE(2) AND ceros_ok(14)) OR (outputF(2) AND ceros_ok(15));
			registro_final(35) <= (output0(3) AND ceros_ok(0)) OR (output1(3) AND ceros_ok(1)) OR (output2(3) AND ceros_ok(2)) OR (output3(3) AND ceros_ok(3)) OR (output4(3) AND ceros_ok(4)) OR (output5(3) AND ceros_ok(5)) OR (output6(3) AND ceros_ok(6)) OR (output7(3) AND ceros_ok(7))OR (output8(3) AND ceros_ok(8))OR (output9(3) AND ceros_ok(9)) OR (outputA(3) AND ceros_ok(10)) OR (outputB(3) AND ceros_ok(11)) OR (outputC(3) AND ceros_ok(12)) OR (outputD(3) AND ceros_ok(13)) OR (outputE(3) AND ceros_ok(14)) OR (outputF(3) AND ceros_ok(15));
			registro_final(36) <= (output0(4) AND ceros_ok(0)) OR (output1(4) AND ceros_ok(1)) OR (output2(4) AND ceros_ok(2)) OR (output3(4) AND ceros_ok(3)) OR (output4(4) AND ceros_ok(4)) OR (output5(4) AND ceros_ok(5)) OR (output6(4) AND ceros_ok(6)) OR (output7(4) AND ceros_ok(7))OR (output8(4) AND ceros_ok(8))OR (output9(4) AND ceros_ok(9)) OR (outputA(4) AND ceros_ok(10)) OR (outputB(4) AND ceros_ok(11)) OR (outputC(4) AND ceros_ok(12)) OR (outputD(4) AND ceros_ok(13)) OR (outputE(4) AND ceros_ok(14)) OR (outputF(4) AND ceros_ok(15));
			registro_final(37) <= (output0(5) AND ceros_ok(0)) OR (output1(5) AND ceros_ok(1)) OR (output2(5) AND ceros_ok(2)) OR (output3(5) AND ceros_ok(3)) OR (output4(5) AND ceros_ok(4)) OR (output5(5) AND ceros_ok(5)) OR (output6(5) AND ceros_ok(6)) OR (output7(5) AND ceros_ok(7))OR (output8(5) AND ceros_ok(8))OR (output9(5) AND ceros_ok(9)) OR (outputA(5) AND ceros_ok(10)) OR (outputB(5) AND ceros_ok(11)) OR (outputC(5) AND ceros_ok(12)) OR (outputD(5) AND ceros_ok(13)) OR (outputE(5) AND ceros_ok(14)) OR (outputF(5) AND ceros_ok(15));
			registro_final(38) <= (output0(6) AND ceros_ok(0)) OR (output1(6) AND ceros_ok(1)) OR (output2(6) AND ceros_ok(2)) OR (output3(6) AND ceros_ok(3)) OR (output4(6) AND ceros_ok(4)) OR (output5(6) AND ceros_ok(5)) OR (output6(6) AND ceros_ok(6)) OR (output7(6) AND ceros_ok(7))OR (output8(6) AND ceros_ok(8))OR (output9(6) AND ceros_ok(9)) OR (outputA(6) AND ceros_ok(10)) OR (outputB(6) AND ceros_ok(11)) OR (outputC(6) AND ceros_ok(12)) OR (outputD(6) AND ceros_ok(13)) OR (outputE(6) AND ceros_ok(14)) OR (outputF(6) AND ceros_ok(15));
			registro_final(39) <= (output0(7) AND ceros_ok(0)) OR (output1(7) AND ceros_ok(1)) OR (output2(7) AND ceros_ok(2)) OR (output3(7) AND ceros_ok(3)) OR (output4(7) AND ceros_ok(4)) OR (output5(7) AND ceros_ok(5)) OR (output6(7) AND ceros_ok(6)) OR (output7(7) AND ceros_ok(7))OR (output8(7) AND ceros_ok(8))OR (output9(7) AND ceros_ok(9)) OR (outputA(7) AND ceros_ok(10)) OR (outputB(7) AND ceros_ok(11)) OR (outputC(7) AND ceros_ok(12)) OR (outputD(7) AND ceros_ok(13)) OR (outputE(7) AND ceros_ok(14)) OR (outputF(7) AND ceros_ok(15));
			registro_final(40) <= (output0(8) AND ceros_ok(0)) OR (output1(8) AND ceros_ok(1)) OR (output2(8) AND ceros_ok(2)) OR (output3(8) AND ceros_ok(3)) OR (output4(8) AND ceros_ok(4)) OR (output5(8) AND ceros_ok(5)) OR (output6(8) AND ceros_ok(6)) OR (output7(8) AND ceros_ok(7))OR (output8(8) AND ceros_ok(8))OR (output9(8) AND ceros_ok(9)) OR (outputA(8) AND ceros_ok(10)) OR (outputB(8) AND ceros_ok(11)) OR (outputC(8) AND ceros_ok(12)) OR (outputD(8) AND ceros_ok(13)) OR (outputE(8) AND ceros_ok(14)) OR (outputF(8) AND ceros_ok(15));
			registro_final(41) <= (output0(9) AND ceros_ok(0)) OR (output1(9) AND ceros_ok(1)) OR (output2(9) AND ceros_ok(2)) OR (output3(9) AND ceros_ok(3)) OR (output4(9) AND ceros_ok(4)) OR (output5(9) AND ceros_ok(5)) OR (output6(9) AND ceros_ok(6)) OR (output7(9) AND ceros_ok(7))OR (output8(9) AND ceros_ok(8))OR (output9(9) AND ceros_ok(9)) OR (outputA(9) AND ceros_ok(10)) OR (outputB(9) AND ceros_ok(11)) OR (outputC(9) AND ceros_ok(12)) OR (outputD(9) AND ceros_ok(13)) OR (outputE(9) AND ceros_ok(14)) OR (outputF(9) AND ceros_ok(15));
			registro_final(42) <= (output0(10) AND ceros_ok(0)) OR (output1(10) AND ceros_ok(1)) OR (output2(10) AND ceros_ok(2)) OR (output3(10) AND ceros_ok(3)) OR (output4(10) AND ceros_ok(4)) OR (output5(10) AND ceros_ok(5)) OR (output6(10) AND ceros_ok(6)) OR (output7(10) AND ceros_ok(7))OR (output8(10) AND ceros_ok(8))OR (output9(10) AND ceros_ok(9)) OR (outputA(10) AND ceros_ok(10)) OR (outputB(10) AND ceros_ok(11)) OR (outputC(10) AND ceros_ok(12)) OR (outputD(10) AND ceros_ok(13)) OR (outputE(10) AND ceros_ok(14)) OR (outputF(10) AND ceros_ok(15));
			registro_final(43) <= (output0(11) AND ceros_ok(0)) OR (output1(11) AND ceros_ok(1)) OR (output2(11) AND ceros_ok(2)) OR (output3(11) AND ceros_ok(3)) OR (output4(11) AND ceros_ok(4)) OR (output5(11) AND ceros_ok(5)) OR (output6(11) AND ceros_ok(6)) OR (output7(11) AND ceros_ok(7))OR (output8(11) AND ceros_ok(8))OR (output9(11) AND ceros_ok(9)) OR (outputA(11) AND ceros_ok(10)) OR (outputB(11) AND ceros_ok(11)) OR (outputC(11) AND ceros_ok(12)) OR (outputD(11) AND ceros_ok(13)) OR (outputE(11) AND ceros_ok(14)) OR (outputF(11) AND ceros_ok(15));
			registro_final(44) <= (output0(12) AND ceros_ok(0)) OR (output1(12) AND ceros_ok(1)) OR (output2(12) AND ceros_ok(2)) OR (output3(12) AND ceros_ok(3)) OR (output4(12) AND ceros_ok(4)) OR (output5(12) AND ceros_ok(5)) OR (output6(12) AND ceros_ok(6)) OR (output7(12) AND ceros_ok(7))OR (output8(12) AND ceros_ok(8))OR (output9(12) AND ceros_ok(9)) OR (outputA(12) AND ceros_ok(10)) OR (outputB(12) AND ceros_ok(11)) OR (outputC(12) AND ceros_ok(12)) OR (outputD(12) AND ceros_ok(13)) OR (outputE(12) AND ceros_ok(14)) OR (outputF(12) AND ceros_ok(15));
			registro_final(45) <= (output0(13) AND ceros_ok(0)) OR (output1(13) AND ceros_ok(1)) OR (output2(13) AND ceros_ok(2)) OR (output3(13) AND ceros_ok(3)) OR (output4(13) AND ceros_ok(4)) OR (output5(13) AND ceros_ok(5)) OR (output6(13) AND ceros_ok(6)) OR (output7(13) AND ceros_ok(7))OR (output8(13) AND ceros_ok(8))OR (output9(13) AND ceros_ok(9)) OR (outputA(13) AND ceros_ok(10)) OR (outputB(13) AND ceros_ok(11)) OR (outputC(13) AND ceros_ok(12)) OR (outputD(13) AND ceros_ok(13)) OR (outputE(13) AND ceros_ok(14)) OR (outputF(13) AND ceros_ok(15));
			registro_final(46) <= (output0(14) AND ceros_ok(0)) OR (output1(14) AND ceros_ok(1)) OR (output2(14) AND ceros_ok(2)) OR (output3(14) AND ceros_ok(3)) OR (output4(14) AND ceros_ok(4)) OR (output5(14) AND ceros_ok(5)) OR (output6(14) AND ceros_ok(6)) OR (output7(14) AND ceros_ok(7))OR (output8(14) AND ceros_ok(8))OR (output9(14) AND ceros_ok(9)) OR (outputA(14) AND ceros_ok(10)) OR (outputB(14) AND ceros_ok(11)) OR (outputC(14) AND ceros_ok(12)) OR (outputD(14) AND ceros_ok(13)) OR (outputE(14) AND ceros_ok(14)) OR (outputF(14) AND ceros_ok(15));
			registro_final(47) <= (output0(15) AND ceros_ok(0)) OR (output1(15) AND ceros_ok(1)) OR (output2(15) AND ceros_ok(2)) OR (output3(15) AND ceros_ok(3)) OR (output4(15) AND ceros_ok(4)) OR (output5(15) AND ceros_ok(5)) OR (output6(15) AND ceros_ok(6)) OR (output7(15) AND ceros_ok(7))OR (output8(15) AND ceros_ok(8))OR (output9(15) AND ceros_ok(9)) OR (outputA(15) AND ceros_ok(10)) OR (outputB(15) AND ceros_ok(11)) OR (outputC(15) AND ceros_ok(12)) OR (outputD(15) AND ceros_ok(13)) OR (outputE(15) AND ceros_ok(14)) OR (outputF(15) AND ceros_ok(15));
			registro_final(48) <= (output0(16) AND ceros_ok(0)) OR (output1(16) AND ceros_ok(1)) OR (output2(16) AND ceros_ok(2)) OR (output3(16) AND ceros_ok(3)) OR (output4(16) AND ceros_ok(4)) OR (output5(16) AND ceros_ok(5)) OR (output6(16) AND ceros_ok(6)) OR (output7(16) AND ceros_ok(7))OR (output8(16) AND ceros_ok(8))OR (output9(16) AND ceros_ok(9)) OR (outputA(16) AND ceros_ok(10)) OR (outputB(16) AND ceros_ok(11)) OR (outputC(16) AND ceros_ok(12)) OR (outputD(16) AND ceros_ok(13)) OR (outputE(16) AND ceros_ok(14)) OR (outputF(16) AND ceros_ok(15));
			registro_final(49) <= (output0(17) AND ceros_ok(0)) OR (output1(17) AND ceros_ok(1)) OR (output2(17) AND ceros_ok(2)) OR (output3(17) AND ceros_ok(3)) OR (output4(17) AND ceros_ok(4)) OR (output5(17) AND ceros_ok(5)) OR (output6(17) AND ceros_ok(6)) OR (output7(17) AND ceros_ok(7))OR (output8(17) AND ceros_ok(8))OR (output9(17) AND ceros_ok(9)) OR (outputA(17) AND ceros_ok(10)) OR (outputB(17) AND ceros_ok(11)) OR (outputC(17) AND ceros_ok(12)) OR (outputD(17) AND ceros_ok(13)) OR (outputE(17) AND ceros_ok(14)) OR (outputF(17) AND ceros_ok(15));
			registro_final(50) <= (output0(18) AND ceros_ok(0)) OR (output1(18) AND ceros_ok(1)) OR (output2(18) AND ceros_ok(2)) OR (output3(18) AND ceros_ok(3)) OR (output4(18) AND ceros_ok(4)) OR (output5(18) AND ceros_ok(5)) OR (output6(18) AND ceros_ok(6)) OR (output7(18) AND ceros_ok(7))OR (output8(18) AND ceros_ok(8))OR (output9(18) AND ceros_ok(9)) OR (outputA(18) AND ceros_ok(10)) OR (outputB(18) AND ceros_ok(11)) OR (outputC(18) AND ceros_ok(12)) OR (outputD(18) AND ceros_ok(13)) OR (outputE(18) AND ceros_ok(14)) OR (outputF(18) AND ceros_ok(15));
			registro_final(51) <= (output0(19) AND ceros_ok(0)) OR (output1(19) AND ceros_ok(1)) OR (output2(19) AND ceros_ok(2)) OR (output3(19) AND ceros_ok(3)) OR (output4(19) AND ceros_ok(4)) OR (output5(19) AND ceros_ok(5)) OR (output6(19) AND ceros_ok(6)) OR (output7(19) AND ceros_ok(7))OR (output8(19) AND ceros_ok(8))OR (output9(19) AND ceros_ok(9)) OR (outputA(19) AND ceros_ok(10)) OR (outputB(19) AND ceros_ok(11)) OR (outputC(19) AND ceros_ok(12)) OR (outputD(19) AND ceros_ok(13)) OR (outputE(19) AND ceros_ok(14)) OR (outputF(19) AND ceros_ok(15));
			registro_final(52) <= (output0(20) AND ceros_ok(0)) OR (output1(20) AND ceros_ok(1)) OR (output2(20) AND ceros_ok(2)) OR (output3(20) AND ceros_ok(3)) OR (output4(20) AND ceros_ok(4)) OR (output5(20) AND ceros_ok(5)) OR (output6(20) AND ceros_ok(6)) OR (output7(20) AND ceros_ok(7))OR (output8(20) AND ceros_ok(8))OR (output9(20) AND ceros_ok(9)) OR (outputA(20) AND ceros_ok(10)) OR (outputB(20) AND ceros_ok(11)) OR (outputC(20) AND ceros_ok(12)) OR (outputD(20) AND ceros_ok(13)) OR (outputE(20) AND ceros_ok(14)) OR (outputF(20) AND ceros_ok(15));
			registro_final(53) <= (output0(21) AND ceros_ok(0)) OR (output1(21) AND ceros_ok(1)) OR (output2(21) AND ceros_ok(2)) OR (output3(21) AND ceros_ok(3)) OR (output4(21) AND ceros_ok(4)) OR (output5(21) AND ceros_ok(5)) OR (output6(21) AND ceros_ok(6)) OR (output7(21) AND ceros_ok(7))OR (output8(21) AND ceros_ok(8))OR (output9(21) AND ceros_ok(9)) OR (outputA(21) AND ceros_ok(10)) OR (outputB(21) AND ceros_ok(11)) OR (outputC(21) AND ceros_ok(12)) OR (outputD(21) AND ceros_ok(13)) OR (outputE(21) AND ceros_ok(14)) OR (outputF(21) AND ceros_ok(15));
			registro_final(54) <= (output0(22) AND ceros_ok(0)) OR (output1(22) AND ceros_ok(1)) OR (output2(22) AND ceros_ok(2)) OR (output3(22) AND ceros_ok(3)) OR (output4(22) AND ceros_ok(4)) OR (output5(22) AND ceros_ok(5)) OR (output6(22) AND ceros_ok(6)) OR (output7(22) AND ceros_ok(7))OR (output8(22) AND ceros_ok(8))OR (output9(22) AND ceros_ok(9)) OR (outputA(22) AND ceros_ok(10)) OR (outputB(22) AND ceros_ok(11)) OR (outputC(22) AND ceros_ok(12)) OR (outputD(22) AND ceros_ok(13)) OR (outputE(22) AND ceros_ok(14)) OR (outputF(22) AND ceros_ok(15));
			registro_final(55) <= (output0(23) AND ceros_ok(0)) OR (output1(23) AND ceros_ok(1)) OR (output2(23) AND ceros_ok(2)) OR (output3(23) AND ceros_ok(3)) OR (output4(23) AND ceros_ok(4)) OR (output5(23) AND ceros_ok(5)) OR (output6(23) AND ceros_ok(6)) OR (output7(23) AND ceros_ok(7))OR (output8(23) AND ceros_ok(8))OR (output9(23) AND ceros_ok(9)) OR (outputA(23) AND ceros_ok(10)) OR (outputB(23) AND ceros_ok(11)) OR (outputC(23) AND ceros_ok(12)) OR (outputD(23) AND ceros_ok(13)) OR (outputE(23) AND ceros_ok(14)) OR (outputF(23) AND ceros_ok(15));
			registro_final(56) <= (output0(24) AND ceros_ok(0)) OR (output1(24) AND ceros_ok(1)) OR (output2(24) AND ceros_ok(2)) OR (output3(24) AND ceros_ok(3)) OR (output4(24) AND ceros_ok(4)) OR (output5(24) AND ceros_ok(5)) OR (output6(24) AND ceros_ok(6)) OR (output7(24) AND ceros_ok(7))OR (output8(24) AND ceros_ok(8))OR (output9(24) AND ceros_ok(9)) OR (outputA(24) AND ceros_ok(10)) OR (outputB(24) AND ceros_ok(11)) OR (outputC(24) AND ceros_ok(12)) OR (outputD(24) AND ceros_ok(13)) OR (outputE(24) AND ceros_ok(14)) OR (outputF(24) AND ceros_ok(15));
			registro_final(57) <= (output0(25) AND ceros_ok(0)) OR (output1(25) AND ceros_ok(1)) OR (output2(25) AND ceros_ok(2)) OR (output3(25) AND ceros_ok(3)) OR (output4(25) AND ceros_ok(4)) OR (output5(25) AND ceros_ok(5)) OR (output6(25) AND ceros_ok(6)) OR (output7(25) AND ceros_ok(7))OR (output8(25) AND ceros_ok(8))OR (output9(25) AND ceros_ok(9)) OR (outputA(25) AND ceros_ok(10)) OR (outputB(25) AND ceros_ok(11)) OR (outputC(25) AND ceros_ok(12)) OR (outputD(25) AND ceros_ok(13)) OR (outputE(25) AND ceros_ok(14)) OR (outputF(25) AND ceros_ok(15));
			registro_final(58) <= (output0(26) AND ceros_ok(0)) OR (output1(26) AND ceros_ok(1)) OR (output2(26) AND ceros_ok(2)) OR (output3(26) AND ceros_ok(3)) OR (output4(26) AND ceros_ok(4)) OR (output5(26) AND ceros_ok(5)) OR (output6(26) AND ceros_ok(6)) OR (output7(26) AND ceros_ok(7))OR (output8(26) AND ceros_ok(8))OR (output9(26) AND ceros_ok(9)) OR (outputA(26) AND ceros_ok(10)) OR (outputB(26) AND ceros_ok(11)) OR (outputC(26) AND ceros_ok(12)) OR (outputD(26) AND ceros_ok(13)) OR (outputE(26) AND ceros_ok(14)) OR (outputF(26) AND ceros_ok(15));
			registro_final(59) <= (output0(27) AND ceros_ok(0)) OR (output1(27) AND ceros_ok(1)) OR (output2(27) AND ceros_ok(2)) OR (output3(27) AND ceros_ok(3)) OR (output4(27) AND ceros_ok(4)) OR (output5(27) AND ceros_ok(5)) OR (output6(27) AND ceros_ok(6)) OR (output7(27) AND ceros_ok(7))OR (output8(27) AND ceros_ok(8))OR (output9(27) AND ceros_ok(9)) OR (outputA(27) AND ceros_ok(10)) OR (outputB(27) AND ceros_ok(11)) OR (outputC(27) AND ceros_ok(12)) OR (outputD(27) AND ceros_ok(13)) OR (outputE(27) AND ceros_ok(14)) OR (outputF(27) AND ceros_ok(15));
			registro_final(60) <= (output0(28) AND ceros_ok(0)) OR (output1(28) AND ceros_ok(1)) OR (output2(28) AND ceros_ok(2)) OR (output3(28) AND ceros_ok(3)) OR (output4(28) AND ceros_ok(4)) OR (output5(28) AND ceros_ok(5)) OR (output6(28) AND ceros_ok(6)) OR (output7(28) AND ceros_ok(7))OR (output8(28) AND ceros_ok(8))OR (output9(28) AND ceros_ok(9)) OR (outputA(28) AND ceros_ok(10)) OR (outputB(28) AND ceros_ok(11)) OR (outputC(28) AND ceros_ok(12)) OR (outputD(28) AND ceros_ok(13)) OR (outputE(28) AND ceros_ok(14)) OR (outputF(28) AND ceros_ok(15));
			registro_final(61) <= (output0(29) AND ceros_ok(0)) OR (output1(29) AND ceros_ok(1)) OR (output2(29) AND ceros_ok(2)) OR (output3(29) AND ceros_ok(3)) OR (output4(29) AND ceros_ok(4)) OR (output5(29) AND ceros_ok(5)) OR (output6(29) AND ceros_ok(6)) OR (output7(29) AND ceros_ok(7))OR (output8(29) AND ceros_ok(8))OR (output9(29) AND ceros_ok(9)) OR (outputA(29) AND ceros_ok(10)) OR (outputB(29) AND ceros_ok(11)) OR (outputC(29) AND ceros_ok(12)) OR (outputD(29) AND ceros_ok(13)) OR (outputE(29) AND ceros_ok(14)) OR (outputF(29) AND ceros_ok(15));
			registro_final(62) <= (output0(30) AND ceros_ok(0)) OR (output1(30) AND ceros_ok(1)) OR (output2(30) AND ceros_ok(2)) OR (output3(30) AND ceros_ok(3)) OR (output4(30) AND ceros_ok(4)) OR (output5(30) AND ceros_ok(5)) OR (output6(30) AND ceros_ok(6)) OR (output7(30) AND ceros_ok(7))OR (output8(30) AND ceros_ok(8))OR (output9(30) AND ceros_ok(9)) OR (outputA(30) AND ceros_ok(10)) OR (outputB(30) AND ceros_ok(11)) OR (outputC(30) AND ceros_ok(12)) OR (outputD(30) AND ceros_ok(13)) OR (outputE(30) AND ceros_ok(14)) OR (outputF(30) AND ceros_ok(15));
			registro_final(63) <= (output0(31) AND ceros_ok(0)) OR (output1(31) AND ceros_ok(1)) OR (output2(31) AND ceros_ok(2)) OR (output3(31) AND ceros_ok(3)) OR (output4(31) AND ceros_ok(4)) OR (output5(31) AND ceros_ok(5)) OR (output6(31) AND ceros_ok(6)) OR (output7(31) AND ceros_ok(7))OR (output8(31) AND ceros_ok(8))OR (output9(31) AND ceros_ok(9)) OR (outputA(31) AND ceros_ok(10)) OR (outputB(31) AND ceros_ok(11)) OR (outputC(31) AND ceros_ok(12)) OR (outputD(31) AND ceros_ok(13)) OR (outputE(31) AND ceros_ok(14)) OR (outputF(31) AND ceros_ok(15));
			registro_final(64) <= (output0(32) AND ceros_ok(0)) OR (output1(32) AND ceros_ok(1)) OR (output2(32) AND ceros_ok(2)) OR (output3(32) AND ceros_ok(3)) OR (output4(32) AND ceros_ok(4)) OR (output5(32) AND ceros_ok(5)) OR (output6(32) AND ceros_ok(6)) OR (output7(32) AND ceros_ok(7))OR (output8(32) AND ceros_ok(8))OR (output9(32) AND ceros_ok(9)) OR (outputA(32) AND ceros_ok(10)) OR (outputB(32) AND ceros_ok(11)) OR (outputC(32) AND ceros_ok(12)) OR (outputD(32) AND ceros_ok(13)) OR (outputE(32) AND ceros_ok(14)) OR (outputF(32) AND ceros_ok(15));
			registro_final(65) <= (output0(33) AND ceros_ok(0)) OR (output1(33) AND ceros_ok(1)) OR (output2(33) AND ceros_ok(2)) OR (output3(33) AND ceros_ok(3)) OR (output4(33) AND ceros_ok(4)) OR (output5(33) AND ceros_ok(5)) OR (output6(33) AND ceros_ok(6)) OR (output7(33) AND ceros_ok(7))OR (output8(33) AND ceros_ok(8))OR (output9(33) AND ceros_ok(9)) OR (outputA(33) AND ceros_ok(10)) OR (outputB(33) AND ceros_ok(11)) OR (outputC(33) AND ceros_ok(12)) OR (outputD(33) AND ceros_ok(13)) OR (outputE(33) AND ceros_ok(14)) OR (outputF(33) AND ceros_ok(15));
			registro_final(66) <= (output0(34) AND ceros_ok(0)) OR (output1(34) AND ceros_ok(1)) OR (output2(34) AND ceros_ok(2)) OR (output3(34) AND ceros_ok(3)) OR (output4(34) AND ceros_ok(4)) OR (output5(34) AND ceros_ok(5)) OR (output6(34) AND ceros_ok(6)) OR (output7(34) AND ceros_ok(7))OR (output8(34) AND ceros_ok(8))OR (output9(34) AND ceros_ok(9)) OR (outputA(34) AND ceros_ok(10)) OR (outputB(34) AND ceros_ok(11)) OR (outputC(34) AND ceros_ok(12)) OR (outputD(34) AND ceros_ok(13)) OR (outputE(34) AND ceros_ok(14)) OR (outputF(34) AND ceros_ok(15));
			registro_final(67) <= (output0(35) AND ceros_ok(0)) OR (output1(35) AND ceros_ok(1)) OR (output2(35) AND ceros_ok(2)) OR (output3(35) AND ceros_ok(3)) OR (output4(35) AND ceros_ok(4)) OR (output5(35) AND ceros_ok(5)) OR (output6(35) AND ceros_ok(6)) OR (output7(35) AND ceros_ok(7))OR (output8(35) AND ceros_ok(8))OR (output9(35) AND ceros_ok(9)) OR (outputA(35) AND ceros_ok(10)) OR (outputB(35) AND ceros_ok(11)) OR (outputC(35) AND ceros_ok(12)) OR (outputD(35) AND ceros_ok(13)) OR (outputE(35) AND ceros_ok(14)) OR (outputF(35) AND ceros_ok(15));
			registro_final(68) <= (output0(36) AND ceros_ok(0)) OR (output1(36) AND ceros_ok(1)) OR (output2(36) AND ceros_ok(2)) OR (output3(36) AND ceros_ok(3)) OR (output4(36) AND ceros_ok(4)) OR (output5(36) AND ceros_ok(5)) OR (output6(36) AND ceros_ok(6)) OR (output7(36) AND ceros_ok(7))OR (output8(36) AND ceros_ok(8))OR (output9(36) AND ceros_ok(9)) OR (outputA(36) AND ceros_ok(10)) OR (outputB(36) AND ceros_ok(11)) OR (outputC(36) AND ceros_ok(12)) OR (outputD(36) AND ceros_ok(13)) OR (outputE(36) AND ceros_ok(14)) OR (outputF(36) AND ceros_ok(15));
			registro_final(69) <= (output0(37) AND ceros_ok(0)) OR (output1(37) AND ceros_ok(1)) OR (output2(37) AND ceros_ok(2)) OR (output3(37) AND ceros_ok(3)) OR (output4(37) AND ceros_ok(4)) OR (output5(37) AND ceros_ok(5)) OR (output6(37) AND ceros_ok(6)) OR (output7(37) AND ceros_ok(7))OR (output8(37) AND ceros_ok(8))OR (output9(37) AND ceros_ok(9)) OR (outputA(37) AND ceros_ok(10)) OR (outputB(37) AND ceros_ok(11)) OR (outputC(37) AND ceros_ok(12)) OR (outputD(37) AND ceros_ok(13)) OR (outputE(37) AND ceros_ok(14)) OR (outputF(37) AND ceros_ok(15));
			registro_final(70) <= (output0(38) AND ceros_ok(0)) OR (output1(38) AND ceros_ok(1)) OR (output2(38) AND ceros_ok(2)) OR (output3(38) AND ceros_ok(3)) OR (output4(38) AND ceros_ok(4)) OR (output5(38) AND ceros_ok(5)) OR (output6(38) AND ceros_ok(6)) OR (output7(38) AND ceros_ok(7))OR (output8(38) AND ceros_ok(8))OR (output9(38) AND ceros_ok(9)) OR (outputA(38) AND ceros_ok(10)) OR (outputB(38) AND ceros_ok(11)) OR (outputC(38) AND ceros_ok(12)) OR (outputD(38) AND ceros_ok(13)) OR (outputE(38) AND ceros_ok(14)) OR (outputF(38) AND ceros_ok(15));
			registro_final(71) <= (output0(39) AND ceros_ok(0)) OR (output1(39) AND ceros_ok(1)) OR (output2(39) AND ceros_ok(2)) OR (output3(39) AND ceros_ok(3)) OR (output4(39) AND ceros_ok(4)) OR (output5(39) AND ceros_ok(5)) OR (output6(39) AND ceros_ok(6)) OR (output7(39) AND ceros_ok(7))OR (output8(39) AND ceros_ok(8))OR (output9(39) AND ceros_ok(9)) OR (outputA(39) AND ceros_ok(10)) OR (outputB(39) AND ceros_ok(11)) OR (outputC(39) AND ceros_ok(12)) OR (outputD(39) AND ceros_ok(13)) OR (outputE(39) AND ceros_ok(14)) OR (outputF(39) AND ceros_ok(15));
			registro_final(72) <= (output0(40) AND ceros_ok(0)) OR (output1(40) AND ceros_ok(1)) OR (output2(40) AND ceros_ok(2)) OR (output3(40) AND ceros_ok(3)) OR (output4(40) AND ceros_ok(4)) OR (output5(40) AND ceros_ok(5)) OR (output6(40) AND ceros_ok(6)) OR (output7(40) AND ceros_ok(7))OR (output8(40) AND ceros_ok(8))OR (output9(40) AND ceros_ok(9)) OR (outputA(40) AND ceros_ok(10)) OR (outputB(40) AND ceros_ok(11)) OR (outputC(40) AND ceros_ok(12)) OR (outputD(40) AND ceros_ok(13)) OR (outputE(40) AND ceros_ok(14)) OR (outputF(40) AND ceros_ok(15));
			registro_final(73) <= (output0(41) AND ceros_ok(0)) OR (output1(41) AND ceros_ok(1)) OR (output2(41) AND ceros_ok(2)) OR (output3(41) AND ceros_ok(3)) OR (output4(41) AND ceros_ok(4)) OR (output5(41) AND ceros_ok(5)) OR (output6(41) AND ceros_ok(6)) OR (output7(41) AND ceros_ok(7))OR (output8(41) AND ceros_ok(8))OR (output9(41) AND ceros_ok(9)) OR (outputA(41) AND ceros_ok(10)) OR (outputB(41) AND ceros_ok(11)) OR (outputC(41) AND ceros_ok(12)) OR (outputD(41) AND ceros_ok(13)) OR (outputE(41) AND ceros_ok(14)) OR (outputF(41) AND ceros_ok(15));
			registro_final(74) <= (output0(42) AND ceros_ok(0)) OR (output1(42) AND ceros_ok(1)) OR (output2(42) AND ceros_ok(2)) OR (output3(42) AND ceros_ok(3)) OR (output4(42) AND ceros_ok(4)) OR (output5(42) AND ceros_ok(5)) OR (output6(42) AND ceros_ok(6)) OR (output7(42) AND ceros_ok(7))OR (output8(42) AND ceros_ok(8))OR (output9(42) AND ceros_ok(9)) OR (outputA(42) AND ceros_ok(10)) OR (outputB(42) AND ceros_ok(11)) OR (outputC(42) AND ceros_ok(12)) OR (outputD(42) AND ceros_ok(13)) OR (outputE(42) AND ceros_ok(14)) OR (outputF(42) AND ceros_ok(15));
			registro_final(75) <= (output0(43) AND ceros_ok(0)) OR (output1(43) AND ceros_ok(1)) OR (output2(43) AND ceros_ok(2)) OR (output3(43) AND ceros_ok(3)) OR (output4(43) AND ceros_ok(4)) OR (output5(43) AND ceros_ok(5)) OR (output6(43) AND ceros_ok(6)) OR (output7(43) AND ceros_ok(7))OR (output8(43) AND ceros_ok(8))OR (output9(43) AND ceros_ok(9)) OR (outputA(43) AND ceros_ok(10)) OR (outputB(43) AND ceros_ok(11)) OR (outputC(43) AND ceros_ok(12)) OR (outputD(43) AND ceros_ok(13)) OR (outputE(43) AND ceros_ok(14)) OR (outputF(43) AND ceros_ok(15));
			registro_final(76) <= (output0(44) AND ceros_ok(0)) OR (output1(44) AND ceros_ok(1)) OR (output2(44) AND ceros_ok(2)) OR (output3(44) AND ceros_ok(3)) OR (output4(44) AND ceros_ok(4)) OR (output5(44) AND ceros_ok(5)) OR (output6(44) AND ceros_ok(6)) OR (output7(44) AND ceros_ok(7))OR (output8(44) AND ceros_ok(8))OR (output9(44) AND ceros_ok(9)) OR (outputA(44) AND ceros_ok(10)) OR (outputB(44) AND ceros_ok(11)) OR (outputC(44) AND ceros_ok(12)) OR (outputD(44) AND ceros_ok(13)) OR (outputE(44) AND ceros_ok(14)) OR (outputF(44) AND ceros_ok(15));
			registro_final(77) <= (output0(45) AND ceros_ok(0)) OR (output1(45) AND ceros_ok(1)) OR (output2(45) AND ceros_ok(2)) OR (output3(45) AND ceros_ok(3)) OR (output4(45) AND ceros_ok(4)) OR (output5(45) AND ceros_ok(5)) OR (output6(45) AND ceros_ok(6)) OR (output7(45) AND ceros_ok(7))OR (output8(45) AND ceros_ok(8))OR (output9(45) AND ceros_ok(9)) OR (outputA(45) AND ceros_ok(10)) OR (outputB(45) AND ceros_ok(11)) OR (outputC(45) AND ceros_ok(12)) OR (outputD(45) AND ceros_ok(13)) OR (outputE(45) AND ceros_ok(14)) OR (outputF(45) AND ceros_ok(15));
			registro_final(78) <= (output0(46) AND ceros_ok(0)) OR (output1(46) AND ceros_ok(1)) OR (output2(46) AND ceros_ok(2)) OR (output3(46) AND ceros_ok(3)) OR (output4(46) AND ceros_ok(4)) OR (output5(46) AND ceros_ok(5)) OR (output6(46) AND ceros_ok(6)) OR (output7(46) AND ceros_ok(7))OR (output8(46) AND ceros_ok(8))OR (output9(46) AND ceros_ok(9)) OR (outputA(46) AND ceros_ok(10)) OR (outputB(46) AND ceros_ok(11)) OR (outputC(46) AND ceros_ok(12)) OR (outputD(46) AND ceros_ok(13)) OR (outputE(46) AND ceros_ok(14)) OR (outputF(46) AND ceros_ok(15));
			registro_final(79) <= (output0(47) AND ceros_ok(0)) OR (output1(47) AND ceros_ok(1)) OR (output2(47) AND ceros_ok(2)) OR (output3(47) AND ceros_ok(3)) OR (output4(47) AND ceros_ok(4)) OR (output5(47) AND ceros_ok(5)) OR (output6(47) AND ceros_ok(6)) OR (output7(47) AND ceros_ok(7))OR (output8(47) AND ceros_ok(8))OR (output9(47) AND ceros_ok(9)) OR (outputA(47) AND ceros_ok(10)) OR (outputB(47) AND ceros_ok(11)) OR (outputC(47) AND ceros_ok(12)) OR (outputD(47) AND ceros_ok(13)) OR (outputE(47) AND ceros_ok(14)) OR (outputF(47) AND ceros_ok(15));
			registro_final(80) <= (output0(48) AND ceros_ok(0)) OR (output1(48) AND ceros_ok(1)) OR (output2(48) AND ceros_ok(2)) OR (output3(48) AND ceros_ok(3)) OR (output4(48) AND ceros_ok(4)) OR (output5(48) AND ceros_ok(5)) OR (output6(48) AND ceros_ok(6)) OR (output7(48) AND ceros_ok(7))OR (output8(48) AND ceros_ok(8))OR (output9(48) AND ceros_ok(9)) OR (outputA(48) AND ceros_ok(10)) OR (outputB(48) AND ceros_ok(11)) OR (outputC(48) AND ceros_ok(12)) OR (outputD(48) AND ceros_ok(13)) OR (outputE(48) AND ceros_ok(14)) OR (outputF(48) AND ceros_ok(15));
			registro_final(81) <= (output0(49) AND ceros_ok(0)) OR (output1(49) AND ceros_ok(1)) OR (output2(49) AND ceros_ok(2)) OR (output3(49) AND ceros_ok(3)) OR (output4(49) AND ceros_ok(4)) OR (output5(49) AND ceros_ok(5)) OR (output6(49) AND ceros_ok(6)) OR (output7(49) AND ceros_ok(7))OR (output8(49) AND ceros_ok(8))OR (output9(49) AND ceros_ok(9)) OR (outputA(49) AND ceros_ok(10)) OR (outputB(49) AND ceros_ok(11)) OR (outputC(49) AND ceros_ok(12)) OR (outputD(49) AND ceros_ok(13)) OR (outputE(49) AND ceros_ok(14)) OR (outputF(49) AND ceros_ok(15));
			registro_final(82) <= (output0(50) AND ceros_ok(0)) OR (output1(50) AND ceros_ok(1)) OR (output2(50) AND ceros_ok(2)) OR (output3(50) AND ceros_ok(3)) OR (output4(50) AND ceros_ok(4)) OR (output5(50) AND ceros_ok(5)) OR (output6(50) AND ceros_ok(6)) OR (output7(50) AND ceros_ok(7))OR (output8(50) AND ceros_ok(8))OR (output9(50) AND ceros_ok(9)) OR (outputA(50) AND ceros_ok(10)) OR (outputB(50) AND ceros_ok(11)) OR (outputC(50) AND ceros_ok(12)) OR (outputD(50) AND ceros_ok(13)) OR (outputE(50) AND ceros_ok(14)) OR (outputF(50) AND ceros_ok(15));
			registro_final(83) <= (output0(51) AND ceros_ok(0)) OR (output1(51) AND ceros_ok(1)) OR (output2(51) AND ceros_ok(2)) OR (output3(51) AND ceros_ok(3)) OR (output4(51) AND ceros_ok(4)) OR (output5(51) AND ceros_ok(5)) OR (output6(51) AND ceros_ok(6)) OR (output7(51) AND ceros_ok(7))OR (output8(51) AND ceros_ok(8))OR (output9(51) AND ceros_ok(9)) OR (outputA(51) AND ceros_ok(10)) OR (outputB(51) AND ceros_ok(11)) OR (outputC(51) AND ceros_ok(12)) OR (outputD(51) AND ceros_ok(13)) OR (outputE(51) AND ceros_ok(14)) OR (outputF(51) AND ceros_ok(15));
			registro_final(84) <= (output0(52) AND ceros_ok(0)) OR (output1(52) AND ceros_ok(1)) OR (output2(52) AND ceros_ok(2)) OR (output3(52) AND ceros_ok(3)) OR (output4(52) AND ceros_ok(4)) OR (output5(52) AND ceros_ok(5)) OR (output6(52) AND ceros_ok(6)) OR (output7(52) AND ceros_ok(7))OR (output8(52) AND ceros_ok(8))OR (output9(52) AND ceros_ok(9)) OR (outputA(52) AND ceros_ok(10)) OR (outputB(52) AND ceros_ok(11)) OR (outputC(52) AND ceros_ok(12)) OR (outputD(52) AND ceros_ok(13)) OR (outputE(52) AND ceros_ok(14)) OR (outputF(52) AND ceros_ok(15));
			registro_final(85) <= (output0(53) AND ceros_ok(0)) OR (output1(53) AND ceros_ok(1)) OR (output2(53) AND ceros_ok(2)) OR (output3(53) AND ceros_ok(3)) OR (output4(53) AND ceros_ok(4)) OR (output5(53) AND ceros_ok(5)) OR (output6(53) AND ceros_ok(6)) OR (output7(53) AND ceros_ok(7))OR (output8(53) AND ceros_ok(8))OR (output9(53) AND ceros_ok(9)) OR (outputA(53) AND ceros_ok(10)) OR (outputB(53) AND ceros_ok(11)) OR (outputC(53) AND ceros_ok(12)) OR (outputD(53) AND ceros_ok(13)) OR (outputE(53) AND ceros_ok(14)) OR (outputF(53) AND ceros_ok(15));
			registro_final(86) <= (output0(54) AND ceros_ok(0)) OR (output1(54) AND ceros_ok(1)) OR (output2(54) AND ceros_ok(2)) OR (output3(54) AND ceros_ok(3)) OR (output4(54) AND ceros_ok(4)) OR (output5(54) AND ceros_ok(5)) OR (output6(54) AND ceros_ok(6)) OR (output7(54) AND ceros_ok(7))OR (output8(54) AND ceros_ok(8))OR (output9(54) AND ceros_ok(9)) OR (outputA(54) AND ceros_ok(10)) OR (outputB(54) AND ceros_ok(11)) OR (outputC(54) AND ceros_ok(12)) OR (outputD(54) AND ceros_ok(13)) OR (outputE(54) AND ceros_ok(14)) OR (outputF(54) AND ceros_ok(15));
			registro_final(87) <= (output0(55) AND ceros_ok(0)) OR (output1(55) AND ceros_ok(1)) OR (output2(55) AND ceros_ok(2)) OR (output3(55) AND ceros_ok(3)) OR (output4(55) AND ceros_ok(4)) OR (output5(55) AND ceros_ok(5)) OR (output6(55) AND ceros_ok(6)) OR (output7(55) AND ceros_ok(7))OR (output8(55) AND ceros_ok(8))OR (output9(55) AND ceros_ok(9)) OR (outputA(55) AND ceros_ok(10)) OR (outputB(55) AND ceros_ok(11)) OR (outputC(55) AND ceros_ok(12)) OR (outputD(55) AND ceros_ok(13)) OR (outputE(55) AND ceros_ok(14)) OR (outputF(55) AND ceros_ok(15));
			registro_final(88) <= (output0(56) AND ceros_ok(0)) OR (output1(56) AND ceros_ok(1)) OR (output2(56) AND ceros_ok(2)) OR (output3(56) AND ceros_ok(3)) OR (output4(56) AND ceros_ok(4)) OR (output5(56) AND ceros_ok(5)) OR (output6(56) AND ceros_ok(6)) OR (output7(56) AND ceros_ok(7))OR (output8(56) AND ceros_ok(8))OR (output9(56) AND ceros_ok(9)) OR (outputA(56) AND ceros_ok(10)) OR (outputB(56) AND ceros_ok(11)) OR (outputC(56) AND ceros_ok(12)) OR (outputD(56) AND ceros_ok(13)) OR (outputE(56) AND ceros_ok(14)) OR (outputF(56) AND ceros_ok(15));
			registro_final(89) <= (output0(57) AND ceros_ok(0)) OR (output1(57) AND ceros_ok(1)) OR (output2(57) AND ceros_ok(2)) OR (output3(57) AND ceros_ok(3)) OR (output4(57) AND ceros_ok(4)) OR (output5(57) AND ceros_ok(5)) OR (output6(57) AND ceros_ok(6)) OR (output7(57) AND ceros_ok(7))OR (output8(57) AND ceros_ok(8))OR (output9(57) AND ceros_ok(9)) OR (outputA(57) AND ceros_ok(10)) OR (outputB(57) AND ceros_ok(11)) OR (outputC(57) AND ceros_ok(12)) OR (outputD(57) AND ceros_ok(13)) OR (outputE(57) AND ceros_ok(14)) OR (outputF(57) AND ceros_ok(15));
			registro_final(90) <= (output0(58) AND ceros_ok(0)) OR (output1(58) AND ceros_ok(1)) OR (output2(58) AND ceros_ok(2)) OR (output3(58) AND ceros_ok(3)) OR (output4(58) AND ceros_ok(4)) OR (output5(58) AND ceros_ok(5)) OR (output6(58) AND ceros_ok(6)) OR (output7(58) AND ceros_ok(7))OR (output8(58) AND ceros_ok(8))OR (output9(58) AND ceros_ok(9)) OR (outputA(58) AND ceros_ok(10)) OR (outputB(58) AND ceros_ok(11)) OR (outputC(58) AND ceros_ok(12)) OR (outputD(58) AND ceros_ok(13)) OR (outputE(58) AND ceros_ok(14)) OR (outputF(58) AND ceros_ok(15));
			registro_final(91) <= (output0(59) AND ceros_ok(0)) OR (output1(59) AND ceros_ok(1)) OR (output2(59) AND ceros_ok(2)) OR (output3(59) AND ceros_ok(3)) OR (output4(59) AND ceros_ok(4)) OR (output5(59) AND ceros_ok(5)) OR (output6(59) AND ceros_ok(6)) OR (output7(59) AND ceros_ok(7))OR (output8(59) AND ceros_ok(8))OR (output9(59) AND ceros_ok(9)) OR (outputA(59) AND ceros_ok(10)) OR (outputB(59) AND ceros_ok(11)) OR (outputC(59) AND ceros_ok(12)) OR (outputD(59) AND ceros_ok(13)) OR (outputE(59) AND ceros_ok(14)) OR (outputF(59) AND ceros_ok(15));
			registro_final(92) <= (output0(60) AND ceros_ok(0)) OR (output1(60) AND ceros_ok(1)) OR (output2(60) AND ceros_ok(2)) OR (output3(60) AND ceros_ok(3)) OR (output4(60) AND ceros_ok(4)) OR (output5(60) AND ceros_ok(5)) OR (output6(60) AND ceros_ok(6)) OR (output7(60) AND ceros_ok(7))OR (output8(60) AND ceros_ok(8))OR (output9(60) AND ceros_ok(9)) OR (outputA(60) AND ceros_ok(10)) OR (outputB(60) AND ceros_ok(11)) OR (outputC(60) AND ceros_ok(12)) OR (outputD(60) AND ceros_ok(13)) OR (outputE(60) AND ceros_ok(14)) OR (outputF(60) AND ceros_ok(15));
			registro_final(93) <= (output0(61) AND ceros_ok(0)) OR (output1(61) AND ceros_ok(1)) OR (output2(61) AND ceros_ok(2)) OR (output3(61) AND ceros_ok(3)) OR (output4(61) AND ceros_ok(4)) OR (output5(61) AND ceros_ok(5)) OR (output6(61) AND ceros_ok(6)) OR (output7(61) AND ceros_ok(7))OR (output8(61) AND ceros_ok(8))OR (output9(61) AND ceros_ok(9)) OR (outputA(61) AND ceros_ok(10)) OR (outputB(61) AND ceros_ok(11)) OR (outputC(61) AND ceros_ok(12)) OR (outputD(61) AND ceros_ok(13)) OR (outputE(61) AND ceros_ok(14)) OR (outputF(61) AND ceros_ok(15));
			registro_final(94) <= (output0(62) AND ceros_ok(0)) OR (output1(62) AND ceros_ok(1)) OR (output2(62) AND ceros_ok(2)) OR (output3(62) AND ceros_ok(3)) OR (output4(62) AND ceros_ok(4)) OR (output5(62) AND ceros_ok(5)) OR (output6(62) AND ceros_ok(6)) OR (output7(62) AND ceros_ok(7))OR (output8(62) AND ceros_ok(8))OR (output9(62) AND ceros_ok(9)) OR (outputA(62) AND ceros_ok(10)) OR (outputB(62) AND ceros_ok(11)) OR (outputC(62) AND ceros_ok(12)) OR (outputD(62) AND ceros_ok(13)) OR (outputE(62) AND ceros_ok(14)) OR (outputF(62) AND ceros_ok(15));
			registro_final(95) <= (output0(63) AND ceros_ok(0)) OR (output1(63) AND ceros_ok(1)) OR (output2(63) AND ceros_ok(2)) OR (output3(63) AND ceros_ok(3)) OR (output4(63) AND ceros_ok(4)) OR (output5(63) AND ceros_ok(5)) OR (output6(63) AND ceros_ok(6)) OR (output7(63) AND ceros_ok(7))OR (output8(63) AND ceros_ok(8))OR (output9(63) AND ceros_ok(9)) OR (outputA(63) AND ceros_ok(10)) OR (outputB(63) AND ceros_ok(11)) OR (outputC(63) AND ceros_ok(12)) OR (outputD(63) AND ceros_ok(13)) OR (outputE(63) AND ceros_ok(14)) OR (outputF(63) AND ceros_ok(15));
			registro_final(96) <= (output0(64) AND ceros_ok(0)) OR (output1(64) AND ceros_ok(1)) OR (output2(64) AND ceros_ok(2)) OR (output3(64) AND ceros_ok(3)) OR (output4(64) AND ceros_ok(4)) OR (output5(64) AND ceros_ok(5)) OR (output6(64) AND ceros_ok(6)) OR (output7(64) AND ceros_ok(7))OR (output8(64) AND ceros_ok(8))OR (output9(64) AND ceros_ok(9)) OR (outputA(64) AND ceros_ok(10)) OR (outputB(64) AND ceros_ok(11)) OR (outputC(64) AND ceros_ok(12)) OR (outputD(64) AND ceros_ok(13)) OR (outputE(64) AND ceros_ok(14)) OR (outputF(64) AND ceros_ok(15));
			registro_final(97) <= (output0(65) AND ceros_ok(0)) OR (output1(65) AND ceros_ok(1)) OR (output2(65) AND ceros_ok(2)) OR (output3(65) AND ceros_ok(3)) OR (output4(65) AND ceros_ok(4)) OR (output5(65) AND ceros_ok(5)) OR (output6(65) AND ceros_ok(6)) OR (output7(65) AND ceros_ok(7))OR (output8(65) AND ceros_ok(8))OR (output9(65) AND ceros_ok(9)) OR (outputA(65) AND ceros_ok(10)) OR (outputB(65) AND ceros_ok(11)) OR (outputC(65) AND ceros_ok(12)) OR (outputD(65) AND ceros_ok(13)) OR (outputE(65) AND ceros_ok(14)) OR (outputF(65) AND ceros_ok(15));
			registro_final(98) <= (output0(66) AND ceros_ok(0)) OR (output1(66) AND ceros_ok(1)) OR (output2(66) AND ceros_ok(2)) OR (output3(66) AND ceros_ok(3)) OR (output4(66) AND ceros_ok(4)) OR (output5(66) AND ceros_ok(5)) OR (output6(66) AND ceros_ok(6)) OR (output7(66) AND ceros_ok(7))OR (output8(66) AND ceros_ok(8))OR (output9(66) AND ceros_ok(9)) OR (outputA(66) AND ceros_ok(10)) OR (outputB(66) AND ceros_ok(11)) OR (outputC(66) AND ceros_ok(12)) OR (outputD(66) AND ceros_ok(13)) OR (outputE(66) AND ceros_ok(14)) OR (outputF(66) AND ceros_ok(15));
			registro_final(99) <= (output0(67) AND ceros_ok(0)) OR (output1(67) AND ceros_ok(1)) OR (output2(67) AND ceros_ok(2)) OR (output3(67) AND ceros_ok(3)) OR (output4(67) AND ceros_ok(4)) OR (output5(67) AND ceros_ok(5)) OR (output6(67) AND ceros_ok(6)) OR (output7(67) AND ceros_ok(7))OR (output8(67) AND ceros_ok(8))OR (output9(67) AND ceros_ok(9)) OR (outputA(67) AND ceros_ok(10)) OR (outputB(67) AND ceros_ok(11)) OR (outputC(67) AND ceros_ok(12)) OR (outputD(67) AND ceros_ok(13)) OR (outputE(67) AND ceros_ok(14)) OR (outputF(67) AND ceros_ok(15));
			registro_final(100) <= (output0(68) AND ceros_ok(0)) OR (output1(68) AND ceros_ok(1)) OR (output2(68) AND ceros_ok(2)) OR (output3(68) AND ceros_ok(3)) OR (output4(68) AND ceros_ok(4)) OR (output5(68) AND ceros_ok(5)) OR (output6(68) AND ceros_ok(6)) OR (output7(68) AND ceros_ok(7))OR (output8(68) AND ceros_ok(8))OR (output9(68) AND ceros_ok(9)) OR (outputA(68) AND ceros_ok(10)) OR (outputB(68) AND ceros_ok(11)) OR (outputC(68) AND ceros_ok(12)) OR (outputD(68) AND ceros_ok(13)) OR (outputE(68) AND ceros_ok(14)) OR (outputF(68) AND ceros_ok(15));
			registro_final(101) <= (output0(69) AND ceros_ok(0)) OR (output1(69) AND ceros_ok(1)) OR (output2(69) AND ceros_ok(2)) OR (output3(69) AND ceros_ok(3)) OR (output4(69) AND ceros_ok(4)) OR (output5(69) AND ceros_ok(5)) OR (output6(69) AND ceros_ok(6)) OR (output7(69) AND ceros_ok(7))OR (output8(69) AND ceros_ok(8))OR (output9(69) AND ceros_ok(9)) OR (outputA(69) AND ceros_ok(10)) OR (outputB(69) AND ceros_ok(11)) OR (outputC(69) AND ceros_ok(12)) OR (outputD(69) AND ceros_ok(13)) OR (outputE(69) AND ceros_ok(14)) OR (outputF(69) AND ceros_ok(15));
			registro_final(102) <= (output0(70) AND ceros_ok(0)) OR (output1(70) AND ceros_ok(1)) OR (output2(70) AND ceros_ok(2)) OR (output3(70) AND ceros_ok(3)) OR (output4(70) AND ceros_ok(4)) OR (output5(70) AND ceros_ok(5)) OR (output6(70) AND ceros_ok(6)) OR (output7(70) AND ceros_ok(7))OR (output8(70) AND ceros_ok(8))OR (output9(70) AND ceros_ok(9)) OR (outputA(70) AND ceros_ok(10)) OR (outputB(70) AND ceros_ok(11)) OR (outputC(70) AND ceros_ok(12)) OR (outputD(70) AND ceros_ok(13)) OR (outputE(70) AND ceros_ok(14)) OR (outputF(70) AND ceros_ok(15));
			registro_final(103) <= (output0(71) AND ceros_ok(0)) OR (output1(71) AND ceros_ok(1)) OR (output2(71) AND ceros_ok(2)) OR (output3(71) AND ceros_ok(3)) OR (output4(71) AND ceros_ok(4)) OR (output5(71) AND ceros_ok(5)) OR (output6(71) AND ceros_ok(6)) OR (output7(71) AND ceros_ok(7))OR (output8(71) AND ceros_ok(8))OR (output9(71) AND ceros_ok(9)) OR (outputA(71) AND ceros_ok(10)) OR (outputB(71) AND ceros_ok(11)) OR (outputC(71) AND ceros_ok(12)) OR (outputD(71) AND ceros_ok(13)) OR (outputE(71) AND ceros_ok(14)) OR (outputF(71) AND ceros_ok(15));
			registro_final(104) <= (output0(72) AND ceros_ok(0)) OR (output1(72) AND ceros_ok(1)) OR (output2(72) AND ceros_ok(2)) OR (output3(72) AND ceros_ok(3)) OR (output4(72) AND ceros_ok(4)) OR (output5(72) AND ceros_ok(5)) OR (output6(72) AND ceros_ok(6)) OR (output7(72) AND ceros_ok(7))OR (output8(72) AND ceros_ok(8))OR (output9(72) AND ceros_ok(9)) OR (outputA(72) AND ceros_ok(10)) OR (outputB(72) AND ceros_ok(11)) OR (outputC(72) AND ceros_ok(12)) OR (outputD(72) AND ceros_ok(13)) OR (outputE(72) AND ceros_ok(14)) OR (outputF(72) AND ceros_ok(15));
			registro_final(105) <= (output0(73) AND ceros_ok(0)) OR (output1(73) AND ceros_ok(1)) OR (output2(73) AND ceros_ok(2)) OR (output3(73) AND ceros_ok(3)) OR (output4(73) AND ceros_ok(4)) OR (output5(73) AND ceros_ok(5)) OR (output6(73) AND ceros_ok(6)) OR (output7(73) AND ceros_ok(7))OR (output8(73) AND ceros_ok(8))OR (output9(73) AND ceros_ok(9)) OR (outputA(73) AND ceros_ok(10)) OR (outputB(73) AND ceros_ok(11)) OR (outputC(73) AND ceros_ok(12)) OR (outputD(73) AND ceros_ok(13)) OR (outputE(73) AND ceros_ok(14)) OR (outputF(73) AND ceros_ok(15));
			registro_final(106) <= (output0(74) AND ceros_ok(0)) OR (output1(74) AND ceros_ok(1)) OR (output2(74) AND ceros_ok(2)) OR (output3(74) AND ceros_ok(3)) OR (output4(74) AND ceros_ok(4)) OR (output5(74) AND ceros_ok(5)) OR (output6(74) AND ceros_ok(6)) OR (output7(74) AND ceros_ok(7))OR (output8(74) AND ceros_ok(8))OR (output9(74) AND ceros_ok(9)) OR (outputA(74) AND ceros_ok(10)) OR (outputB(74) AND ceros_ok(11)) OR (outputC(74) AND ceros_ok(12)) OR (outputD(74) AND ceros_ok(13)) OR (outputE(74) AND ceros_ok(14)) OR (outputF(74) AND ceros_ok(15));
			registro_final(107) <= (output0(75) AND ceros_ok(0)) OR (output1(75) AND ceros_ok(1)) OR (output2(75) AND ceros_ok(2)) OR (output3(75) AND ceros_ok(3)) OR (output4(75) AND ceros_ok(4)) OR (output5(75) AND ceros_ok(5)) OR (output6(75) AND ceros_ok(6)) OR (output7(75) AND ceros_ok(7))OR (output8(75) AND ceros_ok(8))OR (output9(75) AND ceros_ok(9)) OR (outputA(75) AND ceros_ok(10)) OR (outputB(75) AND ceros_ok(11)) OR (outputC(75) AND ceros_ok(12)) OR (outputD(75) AND ceros_ok(13)) OR (outputE(75) AND ceros_ok(14)) OR (outputF(75) AND ceros_ok(15));
			registro_final(108) <= (output0(76) AND ceros_ok(0)) OR (output1(76) AND ceros_ok(1)) OR (output2(76) AND ceros_ok(2)) OR (output3(76) AND ceros_ok(3)) OR (output4(76) AND ceros_ok(4)) OR (output5(76) AND ceros_ok(5)) OR (output6(76) AND ceros_ok(6)) OR (output7(76) AND ceros_ok(7))OR (output8(76) AND ceros_ok(8))OR (output9(76) AND ceros_ok(9)) OR (outputA(76) AND ceros_ok(10)) OR (outputB(76) AND ceros_ok(11)) OR (outputC(76) AND ceros_ok(12)) OR (outputD(76) AND ceros_ok(13)) OR (outputE(76) AND ceros_ok(14)) OR (outputF(76) AND ceros_ok(15));
			registro_final(109) <= (output0(77) AND ceros_ok(0)) OR (output1(77) AND ceros_ok(1)) OR (output2(77) AND ceros_ok(2)) OR (output3(77) AND ceros_ok(3)) OR (output4(77) AND ceros_ok(4)) OR (output5(77) AND ceros_ok(5)) OR (output6(77) AND ceros_ok(6)) OR (output7(77) AND ceros_ok(7))OR (output8(77) AND ceros_ok(8))OR (output9(77) AND ceros_ok(9)) OR (outputA(77) AND ceros_ok(10)) OR (outputB(77) AND ceros_ok(11)) OR (outputC(77) AND ceros_ok(12)) OR (outputD(77) AND ceros_ok(13)) OR (outputE(77) AND ceros_ok(14)) OR (outputF(77) AND ceros_ok(15));
			registro_final(110) <= (output0(78) AND ceros_ok(0)) OR (output1(78) AND ceros_ok(1)) OR (output2(78) AND ceros_ok(2)) OR (output3(78) AND ceros_ok(3)) OR (output4(78) AND ceros_ok(4)) OR (output5(78) AND ceros_ok(5)) OR (output6(78) AND ceros_ok(6)) OR (output7(78) AND ceros_ok(7))OR (output8(78) AND ceros_ok(8))OR (output9(78) AND ceros_ok(9)) OR (outputA(78) AND ceros_ok(10)) OR (outputB(78) AND ceros_ok(11)) OR (outputC(78) AND ceros_ok(12)) OR (outputD(78) AND ceros_ok(13)) OR (outputE(78) AND ceros_ok(14)) OR (outputF(78) AND ceros_ok(15));
			registro_final(111) <= (output0(79) AND ceros_ok(0)) OR (output1(79) AND ceros_ok(1)) OR (output2(79) AND ceros_ok(2)) OR (output3(79) AND ceros_ok(3)) OR (output4(79) AND ceros_ok(4)) OR (output5(79) AND ceros_ok(5)) OR (output6(79) AND ceros_ok(6)) OR (output7(79) AND ceros_ok(7))OR (output8(79) AND ceros_ok(8))OR (output9(79) AND ceros_ok(9)) OR (outputA(79) AND ceros_ok(10)) OR (outputB(79) AND ceros_ok(11)) OR (outputC(79) AND ceros_ok(12)) OR (outputD(79) AND ceros_ok(13)) OR (outputE(79) AND ceros_ok(14)) OR (outputF(79) AND ceros_ok(15));
			registro_final(112) <= (output0(80) AND ceros_ok(0)) OR (output1(80) AND ceros_ok(1)) OR (output2(80) AND ceros_ok(2)) OR (output3(80) AND ceros_ok(3)) OR (output4(80) AND ceros_ok(4)) OR (output5(80) AND ceros_ok(5)) OR (output6(80) AND ceros_ok(6)) OR (output7(80) AND ceros_ok(7))OR (output8(80) AND ceros_ok(8))OR (output9(80) AND ceros_ok(9)) OR (outputA(80) AND ceros_ok(10)) OR (outputB(80) AND ceros_ok(11)) OR (outputC(80) AND ceros_ok(12)) OR (outputD(80) AND ceros_ok(13)) OR (outputE(80) AND ceros_ok(14)) OR (outputF(80) AND ceros_ok(15));
			registro_final(113) <= (output0(81) AND ceros_ok(0)) OR (output1(81) AND ceros_ok(1)) OR (output2(81) AND ceros_ok(2)) OR (output3(81) AND ceros_ok(3)) OR (output4(81) AND ceros_ok(4)) OR (output5(81) AND ceros_ok(5)) OR (output6(81) AND ceros_ok(6)) OR (output7(81) AND ceros_ok(7))OR (output8(81) AND ceros_ok(8))OR (output9(81) AND ceros_ok(9)) OR (outputA(81) AND ceros_ok(10)) OR (outputB(81) AND ceros_ok(11)) OR (outputC(81) AND ceros_ok(12)) OR (outputD(81) AND ceros_ok(13)) OR (outputE(81) AND ceros_ok(14)) OR (outputF(81) AND ceros_ok(15));
			registro_final(114) <= (output0(82) AND ceros_ok(0)) OR (output1(82) AND ceros_ok(1)) OR (output2(82) AND ceros_ok(2)) OR (output3(82) AND ceros_ok(3)) OR (output4(82) AND ceros_ok(4)) OR (output5(82) AND ceros_ok(5)) OR (output6(82) AND ceros_ok(6)) OR (output7(82) AND ceros_ok(7))OR (output8(82) AND ceros_ok(8))OR (output9(82) AND ceros_ok(9)) OR (outputA(82) AND ceros_ok(10)) OR (outputB(82) AND ceros_ok(11)) OR (outputC(82) AND ceros_ok(12)) OR (outputD(82) AND ceros_ok(13)) OR (outputE(82) AND ceros_ok(14)) OR (outputF(82) AND ceros_ok(15));
			registro_final(115) <= (output0(83) AND ceros_ok(0)) OR (output1(83) AND ceros_ok(1)) OR (output2(83) AND ceros_ok(2)) OR (output3(83) AND ceros_ok(3)) OR (output4(83) AND ceros_ok(4)) OR (output5(83) AND ceros_ok(5)) OR (output6(83) AND ceros_ok(6)) OR (output7(83) AND ceros_ok(7))OR (output8(83) AND ceros_ok(8))OR (output9(83) AND ceros_ok(9)) OR (outputA(83) AND ceros_ok(10)) OR (outputB(83) AND ceros_ok(11)) OR (outputC(83) AND ceros_ok(12)) OR (outputD(83) AND ceros_ok(13)) OR (outputE(83) AND ceros_ok(14)) OR (outputF(83) AND ceros_ok(15));
			registro_final(116) <= (output0(84) AND ceros_ok(0)) OR (output1(84) AND ceros_ok(1)) OR (output2(84) AND ceros_ok(2)) OR (output3(84) AND ceros_ok(3)) OR (output4(84) AND ceros_ok(4)) OR (output5(84) AND ceros_ok(5)) OR (output6(84) AND ceros_ok(6)) OR (output7(84) AND ceros_ok(7))OR (output8(84) AND ceros_ok(8))OR (output9(84) AND ceros_ok(9)) OR (outputA(84) AND ceros_ok(10)) OR (outputB(84) AND ceros_ok(11)) OR (outputC(84) AND ceros_ok(12)) OR (outputD(84) AND ceros_ok(13)) OR (outputE(84) AND ceros_ok(14)) OR (outputF(84) AND ceros_ok(15));
			registro_final(117) <= (output0(85) AND ceros_ok(0)) OR (output1(85) AND ceros_ok(1)) OR (output2(85) AND ceros_ok(2)) OR (output3(85) AND ceros_ok(3)) OR (output4(85) AND ceros_ok(4)) OR (output5(85) AND ceros_ok(5)) OR (output6(85) AND ceros_ok(6)) OR (output7(85) AND ceros_ok(7))OR (output8(85) AND ceros_ok(8))OR (output9(85) AND ceros_ok(9)) OR (outputA(85) AND ceros_ok(10)) OR (outputB(85) AND ceros_ok(11)) OR (outputC(85) AND ceros_ok(12)) OR (outputD(85) AND ceros_ok(13)) OR (outputE(85) AND ceros_ok(14)) OR (outputF(85) AND ceros_ok(15));
			registro_final(118) <= (output0(86) AND ceros_ok(0)) OR (output1(86) AND ceros_ok(1)) OR (output2(86) AND ceros_ok(2)) OR (output3(86) AND ceros_ok(3)) OR (output4(86) AND ceros_ok(4)) OR (output5(86) AND ceros_ok(5)) OR (output6(86) AND ceros_ok(6)) OR (output7(86) AND ceros_ok(7))OR (output8(86) AND ceros_ok(8))OR (output9(86) AND ceros_ok(9)) OR (outputA(86) AND ceros_ok(10)) OR (outputB(86) AND ceros_ok(11)) OR (outputC(86) AND ceros_ok(12)) OR (outputD(86) AND ceros_ok(13)) OR (outputE(86) AND ceros_ok(14)) OR (outputF(86) AND ceros_ok(15));
			registro_final(119) <= (output0(87) AND ceros_ok(0)) OR (output1(87) AND ceros_ok(1)) OR (output2(87) AND ceros_ok(2)) OR (output3(87) AND ceros_ok(3)) OR (output4(87) AND ceros_ok(4)) OR (output5(87) AND ceros_ok(5)) OR (output6(87) AND ceros_ok(6)) OR (output7(87) AND ceros_ok(7))OR (output8(87) AND ceros_ok(8))OR (output9(87) AND ceros_ok(9)) OR (outputA(87) AND ceros_ok(10)) OR (outputB(87) AND ceros_ok(11)) OR (outputC(87) AND ceros_ok(12)) OR (outputD(87) AND ceros_ok(13)) OR (outputE(87) AND ceros_ok(14)) OR (outputF(87) AND ceros_ok(15));
			registro_final(120) <= (output0(88) AND ceros_ok(0)) OR (output1(88) AND ceros_ok(1)) OR (output2(88) AND ceros_ok(2)) OR (output3(88) AND ceros_ok(3)) OR (output4(88) AND ceros_ok(4)) OR (output5(88) AND ceros_ok(5)) OR (output6(88) AND ceros_ok(6)) OR (output7(88) AND ceros_ok(7))OR (output8(88) AND ceros_ok(8))OR (output9(88) AND ceros_ok(9)) OR (outputA(88) AND ceros_ok(10)) OR (outputB(88) AND ceros_ok(11)) OR (outputC(88) AND ceros_ok(12)) OR (outputD(88) AND ceros_ok(13)) OR (outputE(88) AND ceros_ok(14)) OR (outputF(88) AND ceros_ok(15));
			registro_final(121) <= (output0(89) AND ceros_ok(0)) OR (output1(89) AND ceros_ok(1)) OR (output2(89) AND ceros_ok(2)) OR (output3(89) AND ceros_ok(3)) OR (output4(89) AND ceros_ok(4)) OR (output5(89) AND ceros_ok(5)) OR (output6(89) AND ceros_ok(6)) OR (output7(89) AND ceros_ok(7))OR (output8(89) AND ceros_ok(8))OR (output9(89) AND ceros_ok(9)) OR (outputA(89) AND ceros_ok(10)) OR (outputB(89) AND ceros_ok(11)) OR (outputC(89) AND ceros_ok(12)) OR (outputD(89) AND ceros_ok(13)) OR (outputE(89) AND ceros_ok(14)) OR (outputF(89) AND ceros_ok(15));
			registro_final(122) <= (output0(90) AND ceros_ok(0)) OR (output1(90) AND ceros_ok(1)) OR (output2(90) AND ceros_ok(2)) OR (output3(90) AND ceros_ok(3)) OR (output4(90) AND ceros_ok(4)) OR (output5(90) AND ceros_ok(5)) OR (output6(90) AND ceros_ok(6)) OR (output7(90) AND ceros_ok(7))OR (output8(90) AND ceros_ok(8))OR (output9(90) AND ceros_ok(9)) OR (outputA(90) AND ceros_ok(10)) OR (outputB(90) AND ceros_ok(11)) OR (outputC(90) AND ceros_ok(12)) OR (outputD(90) AND ceros_ok(13)) OR (outputE(90) AND ceros_ok(14)) OR (outputF(90) AND ceros_ok(15));
			registro_final(123) <= (output0(91) AND ceros_ok(0)) OR (output1(91) AND ceros_ok(1)) OR (output2(91) AND ceros_ok(2)) OR (output3(91) AND ceros_ok(3)) OR (output4(91) AND ceros_ok(4)) OR (output5(91) AND ceros_ok(5)) OR (output6(91) AND ceros_ok(6)) OR (output7(91) AND ceros_ok(7))OR (output8(91) AND ceros_ok(8))OR (output9(91) AND ceros_ok(9)) OR (outputA(91) AND ceros_ok(10)) OR (outputB(91) AND ceros_ok(11)) OR (outputC(91) AND ceros_ok(12)) OR (outputD(91) AND ceros_ok(13)) OR (outputE(91) AND ceros_ok(14)) OR (outputF(91) AND ceros_ok(15));
			registro_final(124) <= (output0(92) AND ceros_ok(0)) OR (output1(92) AND ceros_ok(1)) OR (output2(92) AND ceros_ok(2)) OR (output3(92) AND ceros_ok(3)) OR (output4(92) AND ceros_ok(4)) OR (output5(92) AND ceros_ok(5)) OR (output6(92) AND ceros_ok(6)) OR (output7(92) AND ceros_ok(7))OR (output8(92) AND ceros_ok(8))OR (output9(92) AND ceros_ok(9)) OR (outputA(92) AND ceros_ok(10)) OR (outputB(92) AND ceros_ok(11)) OR (outputC(92) AND ceros_ok(12)) OR (outputD(92) AND ceros_ok(13)) OR (outputE(92) AND ceros_ok(14)) OR (outputF(92) AND ceros_ok(15));
			registro_final(125) <= (output0(93) AND ceros_ok(0)) OR (output1(93) AND ceros_ok(1)) OR (output2(93) AND ceros_ok(2)) OR (output3(93) AND ceros_ok(3)) OR (output4(93) AND ceros_ok(4)) OR (output5(93) AND ceros_ok(5)) OR (output6(93) AND ceros_ok(6)) OR (output7(93) AND ceros_ok(7))OR (output8(93) AND ceros_ok(8))OR (output9(93) AND ceros_ok(9)) OR (outputA(93) AND ceros_ok(10)) OR (outputB(93) AND ceros_ok(11)) OR (outputC(93) AND ceros_ok(12)) OR (outputD(93) AND ceros_ok(13)) OR (outputE(93) AND ceros_ok(14)) OR (outputF(93) AND ceros_ok(15));
			registro_final(126) <= (output0(94) AND ceros_ok(0)) OR (output1(94) AND ceros_ok(1)) OR (output2(94) AND ceros_ok(2)) OR (output3(94) AND ceros_ok(3)) OR (output4(94) AND ceros_ok(4)) OR (output5(94) AND ceros_ok(5)) OR (output6(94) AND ceros_ok(6)) OR (output7(94) AND ceros_ok(7))OR (output8(94) AND ceros_ok(8))OR (output9(94) AND ceros_ok(9)) OR (outputA(94) AND ceros_ok(10)) OR (outputB(94) AND ceros_ok(11)) OR (outputC(94) AND ceros_ok(12)) OR (outputD(94) AND ceros_ok(13)) OR (outputE(94) AND ceros_ok(14)) OR (outputF(94) AND ceros_ok(15));
			registro_final(127) <= (output0(95) AND ceros_ok(0)) OR (output1(95) AND ceros_ok(1)) OR (output2(95) AND ceros_ok(2)) OR (output3(95) AND ceros_ok(3)) OR (output4(95) AND ceros_ok(4)) OR (output5(95) AND ceros_ok(5)) OR (output6(95) AND ceros_ok(6)) OR (output7(95) AND ceros_ok(7))OR (output8(95) AND ceros_ok(8))OR (output9(95) AND ceros_ok(9)) OR (outputA(95) AND ceros_ok(10)) OR (outputB(95) AND ceros_ok(11)) OR (outputC(95) AND ceros_ok(12)) OR (outputD(95) AND ceros_ok(13)) OR (outputE(95) AND ceros_ok(14)) OR (outputF(95) AND ceros_ok(15));
			registro_final(128) <= (output0(96) AND ceros_ok(0)) OR (output1(96) AND ceros_ok(1)) OR (output2(96) AND ceros_ok(2)) OR (output3(96) AND ceros_ok(3)) OR (output4(96) AND ceros_ok(4)) OR (output5(96) AND ceros_ok(5)) OR (output6(96) AND ceros_ok(6)) OR (output7(96) AND ceros_ok(7))OR (output8(96) AND ceros_ok(8))OR (output9(96) AND ceros_ok(9)) OR (outputA(96) AND ceros_ok(10)) OR (outputB(96) AND ceros_ok(11)) OR (outputC(96) AND ceros_ok(12)) OR (outputD(96) AND ceros_ok(13)) OR (outputE(96) AND ceros_ok(14)) OR (outputF(96) AND ceros_ok(15));
			registro_final(129) <= (output0(97) AND ceros_ok(0)) OR (output1(97) AND ceros_ok(1)) OR (output2(97) AND ceros_ok(2)) OR (output3(97) AND ceros_ok(3)) OR (output4(97) AND ceros_ok(4)) OR (output5(97) AND ceros_ok(5)) OR (output6(97) AND ceros_ok(6)) OR (output7(97) AND ceros_ok(7))OR (output8(97) AND ceros_ok(8))OR (output9(97) AND ceros_ok(9)) OR (outputA(97) AND ceros_ok(10)) OR (outputB(97) AND ceros_ok(11)) OR (outputC(97) AND ceros_ok(12)) OR (outputD(97) AND ceros_ok(13)) OR (outputE(97) AND ceros_ok(14)) OR (outputF(97) AND ceros_ok(15));
			registro_final(130) <= (output0(98) AND ceros_ok(0)) OR (output1(98) AND ceros_ok(1)) OR (output2(98) AND ceros_ok(2)) OR (output3(98) AND ceros_ok(3)) OR (output4(98) AND ceros_ok(4)) OR (output5(98) AND ceros_ok(5)) OR (output6(98) AND ceros_ok(6)) OR (output7(98) AND ceros_ok(7))OR (output8(98) AND ceros_ok(8))OR (output9(98) AND ceros_ok(9)) OR (outputA(98) AND ceros_ok(10)) OR (outputB(98) AND ceros_ok(11)) OR (outputC(98) AND ceros_ok(12)) OR (outputD(98) AND ceros_ok(13)) OR (outputE(98) AND ceros_ok(14)) OR (outputF(98) AND ceros_ok(15));
			registro_final(131) <= (output0(99) AND ceros_ok(0)) OR (output1(99) AND ceros_ok(1)) OR (output2(99) AND ceros_ok(2)) OR (output3(99) AND ceros_ok(3)) OR (output4(99) AND ceros_ok(4)) OR (output5(99) AND ceros_ok(5)) OR (output6(99) AND ceros_ok(6)) OR (output7(99) AND ceros_ok(7))OR (output8(99) AND ceros_ok(8))OR (output9(99) AND ceros_ok(9)) OR (outputA(99) AND ceros_ok(10)) OR (outputB(99) AND ceros_ok(11)) OR (outputC(99) AND ceros_ok(12)) OR (outputD(99) AND ceros_ok(13)) OR (outputE(99) AND ceros_ok(14)) OR (outputF(99) AND ceros_ok(15));
			registro_final(132) <= (output0(100) AND ceros_ok(0)) OR (output1(100) AND ceros_ok(1)) OR (output2(100) AND ceros_ok(2)) OR (output3(100) AND ceros_ok(3)) OR (output4(100) AND ceros_ok(4)) OR (output5(100) AND ceros_ok(5)) OR (output6(100) AND ceros_ok(6)) OR (output7(100) AND ceros_ok(7))OR (output8(100) AND ceros_ok(8))OR (output9(100) AND ceros_ok(9)) OR (outputA(100) AND ceros_ok(10)) OR (outputB(100) AND ceros_ok(11)) OR (outputC(100) AND ceros_ok(12)) OR (outputD(100) AND ceros_ok(13)) OR (outputE(100) AND ceros_ok(14)) OR (outputF(100) AND ceros_ok(15));
			registro_final(133) <= (output0(101) AND ceros_ok(0)) OR (output1(101) AND ceros_ok(1)) OR (output2(101) AND ceros_ok(2)) OR (output3(101) AND ceros_ok(3)) OR (output4(101) AND ceros_ok(4)) OR (output5(101) AND ceros_ok(5)) OR (output6(101) AND ceros_ok(6)) OR (output7(101) AND ceros_ok(7))OR (output8(101) AND ceros_ok(8))OR (output9(101) AND ceros_ok(9)) OR (outputA(101) AND ceros_ok(10)) OR (outputB(101) AND ceros_ok(11)) OR (outputC(101) AND ceros_ok(12)) OR (outputD(101) AND ceros_ok(13)) OR (outputE(101) AND ceros_ok(14)) OR (outputF(101) AND ceros_ok(15));
			registro_final(134) <= (output0(102) AND ceros_ok(0)) OR (output1(102) AND ceros_ok(1)) OR (output2(102) AND ceros_ok(2)) OR (output3(102) AND ceros_ok(3)) OR (output4(102) AND ceros_ok(4)) OR (output5(102) AND ceros_ok(5)) OR (output6(102) AND ceros_ok(6)) OR (output7(102) AND ceros_ok(7))OR (output8(102) AND ceros_ok(8))OR (output9(102) AND ceros_ok(9)) OR (outputA(102) AND ceros_ok(10)) OR (outputB(102) AND ceros_ok(11)) OR (outputC(102) AND ceros_ok(12)) OR (outputD(102) AND ceros_ok(13)) OR (outputE(102) AND ceros_ok(14)) OR (outputF(102) AND ceros_ok(15));
			registro_final(135) <= (output0(103) AND ceros_ok(0)) OR (output1(103) AND ceros_ok(1)) OR (output2(103) AND ceros_ok(2)) OR (output3(103) AND ceros_ok(3)) OR (output4(103) AND ceros_ok(4)) OR (output5(103) AND ceros_ok(5)) OR (output6(103) AND ceros_ok(6)) OR (output7(103) AND ceros_ok(7))OR (output8(103) AND ceros_ok(8))OR (output9(103) AND ceros_ok(9)) OR (outputA(103) AND ceros_ok(10)) OR (outputB(103) AND ceros_ok(11)) OR (outputC(103) AND ceros_ok(12)) OR (outputD(103) AND ceros_ok(13)) OR (outputE(103) AND ceros_ok(14)) OR (outputF(103) AND ceros_ok(15));
			registro_final(136) <= (output0(104) AND ceros_ok(0)) OR (output1(104) AND ceros_ok(1)) OR (output2(104) AND ceros_ok(2)) OR (output3(104) AND ceros_ok(3)) OR (output4(104) AND ceros_ok(4)) OR (output5(104) AND ceros_ok(5)) OR (output6(104) AND ceros_ok(6)) OR (output7(104) AND ceros_ok(7))OR (output8(104) AND ceros_ok(8))OR (output9(104) AND ceros_ok(9)) OR (outputA(104) AND ceros_ok(10)) OR (outputB(104) AND ceros_ok(11)) OR (outputC(104) AND ceros_ok(12)) OR (outputD(104) AND ceros_ok(13)) OR (outputE(104) AND ceros_ok(14)) OR (outputF(104) AND ceros_ok(15));
			registro_final(137) <= (output0(105) AND ceros_ok(0)) OR (output1(105) AND ceros_ok(1)) OR (output2(105) AND ceros_ok(2)) OR (output3(105) AND ceros_ok(3)) OR (output4(105) AND ceros_ok(4)) OR (output5(105) AND ceros_ok(5)) OR (output6(105) AND ceros_ok(6)) OR (output7(105) AND ceros_ok(7))OR (output8(105) AND ceros_ok(8))OR (output9(105) AND ceros_ok(9)) OR (outputA(105) AND ceros_ok(10)) OR (outputB(105) AND ceros_ok(11)) OR (outputC(105) AND ceros_ok(12)) OR (outputD(105) AND ceros_ok(13)) OR (outputE(105) AND ceros_ok(14)) OR (outputF(105) AND ceros_ok(15));
			registro_final(138) <= (output0(106) AND ceros_ok(0)) OR (output1(106) AND ceros_ok(1)) OR (output2(106) AND ceros_ok(2)) OR (output3(106) AND ceros_ok(3)) OR (output4(106) AND ceros_ok(4)) OR (output5(106) AND ceros_ok(5)) OR (output6(106) AND ceros_ok(6)) OR (output7(106) AND ceros_ok(7))OR (output8(106) AND ceros_ok(8))OR (output9(106) AND ceros_ok(9)) OR (outputA(106) AND ceros_ok(10)) OR (outputB(106) AND ceros_ok(11)) OR (outputC(106) AND ceros_ok(12)) OR (outputD(106) AND ceros_ok(13)) OR (outputE(106) AND ceros_ok(14)) OR (outputF(106) AND ceros_ok(15));
			registro_final(139) <= (output0(107) AND ceros_ok(0)) OR (output1(107) AND ceros_ok(1)) OR (output2(107) AND ceros_ok(2)) OR (output3(107) AND ceros_ok(3)) OR (output4(107) AND ceros_ok(4)) OR (output5(107) AND ceros_ok(5)) OR (output6(107) AND ceros_ok(6)) OR (output7(107) AND ceros_ok(7))OR (output8(107) AND ceros_ok(8))OR (output9(107) AND ceros_ok(9)) OR (outputA(107) AND ceros_ok(10)) OR (outputB(107) AND ceros_ok(11)) OR (outputC(107) AND ceros_ok(12)) OR (outputD(107) AND ceros_ok(13)) OR (outputE(107) AND ceros_ok(14)) OR (outputF(107) AND ceros_ok(15));
			registro_final(140) <= (output0(108) AND ceros_ok(0)) OR (output1(108) AND ceros_ok(1)) OR (output2(108) AND ceros_ok(2)) OR (output3(108) AND ceros_ok(3)) OR (output4(108) AND ceros_ok(4)) OR (output5(108) AND ceros_ok(5)) OR (output6(108) AND ceros_ok(6)) OR (output7(108) AND ceros_ok(7))OR (output8(108) AND ceros_ok(8))OR (output9(108) AND ceros_ok(9)) OR (outputA(108) AND ceros_ok(10)) OR (outputB(108) AND ceros_ok(11)) OR (outputC(108) AND ceros_ok(12)) OR (outputD(108) AND ceros_ok(13)) OR (outputE(108) AND ceros_ok(14)) OR (outputF(108) AND ceros_ok(15));
			registro_final(141) <= (output0(109) AND ceros_ok(0)) OR (output1(109) AND ceros_ok(1)) OR (output2(109) AND ceros_ok(2)) OR (output3(109) AND ceros_ok(3)) OR (output4(109) AND ceros_ok(4)) OR (output5(109) AND ceros_ok(5)) OR (output6(109) AND ceros_ok(6)) OR (output7(109) AND ceros_ok(7))OR (output8(109) AND ceros_ok(8))OR (output9(109) AND ceros_ok(9)) OR (outputA(109) AND ceros_ok(10)) OR (outputB(109) AND ceros_ok(11)) OR (outputC(109) AND ceros_ok(12)) OR (outputD(109) AND ceros_ok(13)) OR (outputE(109) AND ceros_ok(14)) OR (outputF(109) AND ceros_ok(15));
			registro_final(142) <= (output0(110) AND ceros_ok(0)) OR (output1(110) AND ceros_ok(1)) OR (output2(110) AND ceros_ok(2)) OR (output3(110) AND ceros_ok(3)) OR (output4(110) AND ceros_ok(4)) OR (output5(110) AND ceros_ok(5)) OR (output6(110) AND ceros_ok(6)) OR (output7(110) AND ceros_ok(7))OR (output8(110) AND ceros_ok(8))OR (output9(110) AND ceros_ok(9)) OR (outputA(110) AND ceros_ok(10)) OR (outputB(110) AND ceros_ok(11)) OR (outputC(110) AND ceros_ok(12)) OR (outputD(110) AND ceros_ok(13)) OR (outputE(110) AND ceros_ok(14)) OR (outputF(110) AND ceros_ok(15));
			registro_final(143) <= (output0(111) AND ceros_ok(0)) OR (output1(111) AND ceros_ok(1)) OR (output2(111) AND ceros_ok(2)) OR (output3(111) AND ceros_ok(3)) OR (output4(111) AND ceros_ok(4)) OR (output5(111) AND ceros_ok(5)) OR (output6(111) AND ceros_ok(6)) OR (output7(111) AND ceros_ok(7))OR (output8(111) AND ceros_ok(8))OR (output9(111) AND ceros_ok(9)) OR (outputA(111) AND ceros_ok(10)) OR (outputB(111) AND ceros_ok(11)) OR (outputC(111) AND ceros_ok(12)) OR (outputD(111) AND ceros_ok(13)) OR (outputE(111) AND ceros_ok(14)) OR (outputF(111) AND ceros_ok(15));
			registro_final(144) <= (output0(112) AND ceros_ok(0)) OR (output1(112) AND ceros_ok(1)) OR (output2(112) AND ceros_ok(2)) OR (output3(112) AND ceros_ok(3)) OR (output4(112) AND ceros_ok(4)) OR (output5(112) AND ceros_ok(5)) OR (output6(112) AND ceros_ok(6)) OR (output7(112) AND ceros_ok(7))OR (output8(112) AND ceros_ok(8))OR (output9(112) AND ceros_ok(9)) OR (outputA(112) AND ceros_ok(10)) OR (outputB(112) AND ceros_ok(11)) OR (outputC(112) AND ceros_ok(12)) OR (outputD(112) AND ceros_ok(13)) OR (outputE(112) AND ceros_ok(14)) OR (outputF(112) AND ceros_ok(15));
			registro_final(145) <= (output0(113) AND ceros_ok(0)) OR (output1(113) AND ceros_ok(1)) OR (output2(113) AND ceros_ok(2)) OR (output3(113) AND ceros_ok(3)) OR (output4(113) AND ceros_ok(4)) OR (output5(113) AND ceros_ok(5)) OR (output6(113) AND ceros_ok(6)) OR (output7(113) AND ceros_ok(7))OR (output8(113) AND ceros_ok(8))OR (output9(113) AND ceros_ok(9)) OR (outputA(113) AND ceros_ok(10)) OR (outputB(113) AND ceros_ok(11)) OR (outputC(113) AND ceros_ok(12)) OR (outputD(113) AND ceros_ok(13)) OR (outputE(113) AND ceros_ok(14)) OR (outputF(113) AND ceros_ok(15));
			registro_final(146) <= (output0(114) AND ceros_ok(0)) OR (output1(114) AND ceros_ok(1)) OR (output2(114) AND ceros_ok(2)) OR (output3(114) AND ceros_ok(3)) OR (output4(114) AND ceros_ok(4)) OR (output5(114) AND ceros_ok(5)) OR (output6(114) AND ceros_ok(6)) OR (output7(114) AND ceros_ok(7))OR (output8(114) AND ceros_ok(8))OR (output9(114) AND ceros_ok(9)) OR (outputA(114) AND ceros_ok(10)) OR (outputB(114) AND ceros_ok(11)) OR (outputC(114) AND ceros_ok(12)) OR (outputD(114) AND ceros_ok(13)) OR (outputE(114) AND ceros_ok(14)) OR (outputF(114) AND ceros_ok(15));
			registro_final(147) <= (output0(115) AND ceros_ok(0)) OR (output1(115) AND ceros_ok(1)) OR (output2(115) AND ceros_ok(2)) OR (output3(115) AND ceros_ok(3)) OR (output4(115) AND ceros_ok(4)) OR (output5(115) AND ceros_ok(5)) OR (output6(115) AND ceros_ok(6)) OR (output7(115) AND ceros_ok(7))OR (output8(115) AND ceros_ok(8))OR (output9(115) AND ceros_ok(9)) OR (outputA(115) AND ceros_ok(10)) OR (outputB(115) AND ceros_ok(11)) OR (outputC(115) AND ceros_ok(12)) OR (outputD(115) AND ceros_ok(13)) OR (outputE(115) AND ceros_ok(14)) OR (outputF(115) AND ceros_ok(15));
			registro_final(148) <= (output0(116) AND ceros_ok(0)) OR (output1(116) AND ceros_ok(1)) OR (output2(116) AND ceros_ok(2)) OR (output3(116) AND ceros_ok(3)) OR (output4(116) AND ceros_ok(4)) OR (output5(116) AND ceros_ok(5)) OR (output6(116) AND ceros_ok(6)) OR (output7(116) AND ceros_ok(7))OR (output8(116) AND ceros_ok(8))OR (output9(116) AND ceros_ok(9)) OR (outputA(116) AND ceros_ok(10)) OR (outputB(116) AND ceros_ok(11)) OR (outputC(116) AND ceros_ok(12)) OR (outputD(116) AND ceros_ok(13)) OR (outputE(116) AND ceros_ok(14)) OR (outputF(116) AND ceros_ok(15));
			registro_final(149) <= (output0(117) AND ceros_ok(0)) OR (output1(117) AND ceros_ok(1)) OR (output2(117) AND ceros_ok(2)) OR (output3(117) AND ceros_ok(3)) OR (output4(117) AND ceros_ok(4)) OR (output5(117) AND ceros_ok(5)) OR (output6(117) AND ceros_ok(6)) OR (output7(117) AND ceros_ok(7))OR (output8(117) AND ceros_ok(8))OR (output9(117) AND ceros_ok(9)) OR (outputA(117) AND ceros_ok(10)) OR (outputB(117) AND ceros_ok(11)) OR (outputC(117) AND ceros_ok(12)) OR (outputD(117) AND ceros_ok(13)) OR (outputE(117) AND ceros_ok(14)) OR (outputF(117) AND ceros_ok(15));
			registro_final(150) <= (output0(118) AND ceros_ok(0)) OR (output1(118) AND ceros_ok(1)) OR (output2(118) AND ceros_ok(2)) OR (output3(118) AND ceros_ok(3)) OR (output4(118) AND ceros_ok(4)) OR (output5(118) AND ceros_ok(5)) OR (output6(118) AND ceros_ok(6)) OR (output7(118) AND ceros_ok(7))OR (output8(118) AND ceros_ok(8))OR (output9(118) AND ceros_ok(9)) OR (outputA(118) AND ceros_ok(10)) OR (outputB(118) AND ceros_ok(11)) OR (outputC(118) AND ceros_ok(12)) OR (outputD(118) AND ceros_ok(13)) OR (outputE(118) AND ceros_ok(14)) OR (outputF(118) AND ceros_ok(15));
			registro_final(151) <= (output0(119) AND ceros_ok(0)) OR (output1(119) AND ceros_ok(1)) OR (output2(119) AND ceros_ok(2)) OR (output3(119) AND ceros_ok(3)) OR (output4(119) AND ceros_ok(4)) OR (output5(119) AND ceros_ok(5)) OR (output6(119) AND ceros_ok(6)) OR (output7(119) AND ceros_ok(7))OR (output8(119) AND ceros_ok(8))OR (output9(119) AND ceros_ok(9)) OR (outputA(119) AND ceros_ok(10)) OR (outputB(119) AND ceros_ok(11)) OR (outputC(119) AND ceros_ok(12)) OR (outputD(119) AND ceros_ok(13)) OR (outputE(119) AND ceros_ok(14)) OR (outputF(119) AND ceros_ok(15));
			registro_final(152) <= (output0(120) AND ceros_ok(0)) OR (output1(120) AND ceros_ok(1)) OR (output2(120) AND ceros_ok(2)) OR (output3(120) AND ceros_ok(3)) OR (output4(120) AND ceros_ok(4)) OR (output5(120) AND ceros_ok(5)) OR (output6(120) AND ceros_ok(6)) OR (output7(120) AND ceros_ok(7))OR (output8(120) AND ceros_ok(8))OR (output9(120) AND ceros_ok(9)) OR (outputA(120) AND ceros_ok(10)) OR (outputB(120) AND ceros_ok(11)) OR (outputC(120) AND ceros_ok(12)) OR (outputD(120) AND ceros_ok(13)) OR (outputE(120) AND ceros_ok(14)) OR (outputF(120) AND ceros_ok(15));
			registro_final(153) <= (output0(121) AND ceros_ok(0)) OR (output1(121) AND ceros_ok(1)) OR (output2(121) AND ceros_ok(2)) OR (output3(121) AND ceros_ok(3)) OR (output4(121) AND ceros_ok(4)) OR (output5(121) AND ceros_ok(5)) OR (output6(121) AND ceros_ok(6)) OR (output7(121) AND ceros_ok(7))OR (output8(121) AND ceros_ok(8))OR (output9(121) AND ceros_ok(9)) OR (outputA(121) AND ceros_ok(10)) OR (outputB(121) AND ceros_ok(11)) OR (outputC(121) AND ceros_ok(12)) OR (outputD(121) AND ceros_ok(13)) OR (outputE(121) AND ceros_ok(14)) OR (outputF(121) AND ceros_ok(15));
			registro_final(154) <= (output0(122) AND ceros_ok(0)) OR (output1(122) AND ceros_ok(1)) OR (output2(122) AND ceros_ok(2)) OR (output3(122) AND ceros_ok(3)) OR (output4(122) AND ceros_ok(4)) OR (output5(122) AND ceros_ok(5)) OR (output6(122) AND ceros_ok(6)) OR (output7(122) AND ceros_ok(7))OR (output8(122) AND ceros_ok(8))OR (output9(122) AND ceros_ok(9)) OR (outputA(122) AND ceros_ok(10)) OR (outputB(122) AND ceros_ok(11)) OR (outputC(122) AND ceros_ok(12)) OR (outputD(122) AND ceros_ok(13)) OR (outputE(122) AND ceros_ok(14)) OR (outputF(122) AND ceros_ok(15));
			registro_final(155) <= (output0(123) AND ceros_ok(0)) OR (output1(123) AND ceros_ok(1)) OR (output2(123) AND ceros_ok(2)) OR (output3(123) AND ceros_ok(3)) OR (output4(123) AND ceros_ok(4)) OR (output5(123) AND ceros_ok(5)) OR (output6(123) AND ceros_ok(6)) OR (output7(123) AND ceros_ok(7))OR (output8(123) AND ceros_ok(8))OR (output9(123) AND ceros_ok(9)) OR (outputA(123) AND ceros_ok(10)) OR (outputB(123) AND ceros_ok(11)) OR (outputC(123) AND ceros_ok(12)) OR (outputD(123) AND ceros_ok(13)) OR (outputE(123) AND ceros_ok(14)) OR (outputF(123) AND ceros_ok(15));
			registro_final(156) <= (output0(124) AND ceros_ok(0)) OR (output1(124) AND ceros_ok(1)) OR (output2(124) AND ceros_ok(2)) OR (output3(124) AND ceros_ok(3)) OR (output4(124) AND ceros_ok(4)) OR (output5(124) AND ceros_ok(5)) OR (output6(124) AND ceros_ok(6)) OR (output7(124) AND ceros_ok(7))OR (output8(124) AND ceros_ok(8))OR (output9(124) AND ceros_ok(9)) OR (outputA(124) AND ceros_ok(10)) OR (outputB(124) AND ceros_ok(11)) OR (outputC(124) AND ceros_ok(12)) OR (outputD(124) AND ceros_ok(13)) OR (outputE(124) AND ceros_ok(14)) OR (outputF(124) AND ceros_ok(15));
			registro_final(157) <= (output0(125) AND ceros_ok(0)) OR (output1(125) AND ceros_ok(1)) OR (output2(125) AND ceros_ok(2)) OR (output3(125) AND ceros_ok(3)) OR (output4(125) AND ceros_ok(4)) OR (output5(125) AND ceros_ok(5)) OR (output6(125) AND ceros_ok(6)) OR (output7(125) AND ceros_ok(7))OR (output8(125) AND ceros_ok(8))OR (output9(125) AND ceros_ok(9)) OR (outputA(125) AND ceros_ok(10)) OR (outputB(125) AND ceros_ok(11)) OR (outputC(125) AND ceros_ok(12)) OR (outputD(125) AND ceros_ok(13)) OR (outputE(125) AND ceros_ok(14)) OR (outputF(125) AND ceros_ok(15));
			registro_final(158) <= (output0(126) AND ceros_ok(0)) OR (output1(126) AND ceros_ok(1)) OR (output2(126) AND ceros_ok(2)) OR (output3(126) AND ceros_ok(3)) OR (output4(126) AND ceros_ok(4)) OR (output5(126) AND ceros_ok(5)) OR (output6(126) AND ceros_ok(6)) OR (output7(126) AND ceros_ok(7))OR (output8(126) AND ceros_ok(8))OR (output9(126) AND ceros_ok(9)) OR (outputA(126) AND ceros_ok(10)) OR (outputB(126) AND ceros_ok(11)) OR (outputC(126) AND ceros_ok(12)) OR (outputD(126) AND ceros_ok(13)) OR (outputE(126) AND ceros_ok(14)) OR (outputF(126) AND ceros_ok(15));
			registro_final(159) <= (output0(127) AND ceros_ok(0)) OR (output1(127) AND ceros_ok(1)) OR (output2(127) AND ceros_ok(2)) OR (output3(127) AND ceros_ok(3)) OR (output4(127) AND ceros_ok(4)) OR (output5(127) AND ceros_ok(5)) OR (output6(127) AND ceros_ok(6)) OR (output7(127) AND ceros_ok(7))OR (output8(127) AND ceros_ok(8))OR (output9(127) AND ceros_ok(9)) OR (outputA(127) AND ceros_ok(10)) OR (outputB(127) AND ceros_ok(11)) OR (outputC(127) AND ceros_ok(12)) OR (outputD(127) AND ceros_ok(13)) OR (outputE(127) AND ceros_ok(14)) OR (outputF(127) AND ceros_ok(15));
			registro_final(160) <= (output0(128) AND ceros_ok(0)) OR (output1(128) AND ceros_ok(1)) OR (output2(128) AND ceros_ok(2)) OR (output3(128) AND ceros_ok(3)) OR (output4(128) AND ceros_ok(4)) OR (output5(128) AND ceros_ok(5)) OR (output6(128) AND ceros_ok(6)) OR (output7(128) AND ceros_ok(7))OR (output8(128) AND ceros_ok(8))OR (output9(128) AND ceros_ok(9)) OR (outputA(128) AND ceros_ok(10)) OR (outputB(128) AND ceros_ok(11)) OR (outputC(128) AND ceros_ok(12)) OR (outputD(128) AND ceros_ok(13)) OR (outputE(128) AND ceros_ok(14)) OR (outputF(128) AND ceros_ok(15));
			registro_final(161) <= (output0(129) AND ceros_ok(0)) OR (output1(129) AND ceros_ok(1)) OR (output2(129) AND ceros_ok(2)) OR (output3(129) AND ceros_ok(3)) OR (output4(129) AND ceros_ok(4)) OR (output5(129) AND ceros_ok(5)) OR (output6(129) AND ceros_ok(6)) OR (output7(129) AND ceros_ok(7))OR (output8(129) AND ceros_ok(8))OR (output9(129) AND ceros_ok(9)) OR (outputA(129) AND ceros_ok(10)) OR (outputB(129) AND ceros_ok(11)) OR (outputC(129) AND ceros_ok(12)) OR (outputD(129) AND ceros_ok(13)) OR (outputE(129) AND ceros_ok(14)) OR (outputF(129) AND ceros_ok(15));
			registro_final(162) <= (output0(130) AND ceros_ok(0)) OR (output1(130) AND ceros_ok(1)) OR (output2(130) AND ceros_ok(2)) OR (output3(130) AND ceros_ok(3)) OR (output4(130) AND ceros_ok(4)) OR (output5(130) AND ceros_ok(5)) OR (output6(130) AND ceros_ok(6)) OR (output7(130) AND ceros_ok(7))OR (output8(130) AND ceros_ok(8))OR (output9(130) AND ceros_ok(9)) OR (outputA(130) AND ceros_ok(10)) OR (outputB(130) AND ceros_ok(11)) OR (outputC(130) AND ceros_ok(12)) OR (outputD(130) AND ceros_ok(13)) OR (outputE(130) AND ceros_ok(14)) OR (outputF(130) AND ceros_ok(15));
			registro_final(163) <= (output0(131) AND ceros_ok(0)) OR (output1(131) AND ceros_ok(1)) OR (output2(131) AND ceros_ok(2)) OR (output3(131) AND ceros_ok(3)) OR (output4(131) AND ceros_ok(4)) OR (output5(131) AND ceros_ok(5)) OR (output6(131) AND ceros_ok(6)) OR (output7(131) AND ceros_ok(7))OR (output8(131) AND ceros_ok(8))OR (output9(131) AND ceros_ok(9)) OR (outputA(131) AND ceros_ok(10)) OR (outputB(131) AND ceros_ok(11)) OR (outputC(131) AND ceros_ok(12)) OR (outputD(131) AND ceros_ok(13)) OR (outputE(131) AND ceros_ok(14)) OR (outputF(131) AND ceros_ok(15));
			registro_final(164) <= (output0(132) AND ceros_ok(0)) OR (output1(132) AND ceros_ok(1)) OR (output2(132) AND ceros_ok(2)) OR (output3(132) AND ceros_ok(3)) OR (output4(132) AND ceros_ok(4)) OR (output5(132) AND ceros_ok(5)) OR (output6(132) AND ceros_ok(6)) OR (output7(132) AND ceros_ok(7))OR (output8(132) AND ceros_ok(8))OR (output9(132) AND ceros_ok(9)) OR (outputA(132) AND ceros_ok(10)) OR (outputB(132) AND ceros_ok(11)) OR (outputC(132) AND ceros_ok(12)) OR (outputD(132) AND ceros_ok(13)) OR (outputE(132) AND ceros_ok(14)) OR (outputF(132) AND ceros_ok(15));
			registro_final(165) <= (output0(133) AND ceros_ok(0)) OR (output1(133) AND ceros_ok(1)) OR (output2(133) AND ceros_ok(2)) OR (output3(133) AND ceros_ok(3)) OR (output4(133) AND ceros_ok(4)) OR (output5(133) AND ceros_ok(5)) OR (output6(133) AND ceros_ok(6)) OR (output7(133) AND ceros_ok(7))OR (output8(133) AND ceros_ok(8))OR (output9(133) AND ceros_ok(9)) OR (outputA(133) AND ceros_ok(10)) OR (outputB(133) AND ceros_ok(11)) OR (outputC(133) AND ceros_ok(12)) OR (outputD(133) AND ceros_ok(13)) OR (outputE(133) AND ceros_ok(14)) OR (outputF(133) AND ceros_ok(15));
			registro_final(166) <= (output0(134) AND ceros_ok(0)) OR (output1(134) AND ceros_ok(1)) OR (output2(134) AND ceros_ok(2)) OR (output3(134) AND ceros_ok(3)) OR (output4(134) AND ceros_ok(4)) OR (output5(134) AND ceros_ok(5)) OR (output6(134) AND ceros_ok(6)) OR (output7(134) AND ceros_ok(7))OR (output8(134) AND ceros_ok(8))OR (output9(134) AND ceros_ok(9)) OR (outputA(134) AND ceros_ok(10)) OR (outputB(134) AND ceros_ok(11)) OR (outputC(134) AND ceros_ok(12)) OR (outputD(134) AND ceros_ok(13)) OR (outputE(134) AND ceros_ok(14)) OR (outputF(134) AND ceros_ok(15));
			registro_final(167) <= (output0(135) AND ceros_ok(0)) OR (output1(135) AND ceros_ok(1)) OR (output2(135) AND ceros_ok(2)) OR (output3(135) AND ceros_ok(3)) OR (output4(135) AND ceros_ok(4)) OR (output5(135) AND ceros_ok(5)) OR (output6(135) AND ceros_ok(6)) OR (output7(135) AND ceros_ok(7))OR (output8(135) AND ceros_ok(8))OR (output9(135) AND ceros_ok(9)) OR (outputA(135) AND ceros_ok(10)) OR (outputB(135) AND ceros_ok(11)) OR (outputC(135) AND ceros_ok(12)) OR (outputD(135) AND ceros_ok(13)) OR (outputE(135) AND ceros_ok(14)) OR (outputF(135) AND ceros_ok(15));
			registro_final(168) <= (output0(136) AND ceros_ok(0)) OR (output1(136) AND ceros_ok(1)) OR (output2(136) AND ceros_ok(2)) OR (output3(136) AND ceros_ok(3)) OR (output4(136) AND ceros_ok(4)) OR (output5(136) AND ceros_ok(5)) OR (output6(136) AND ceros_ok(6)) OR (output7(136) AND ceros_ok(7))OR (output8(136) AND ceros_ok(8))OR (output9(136) AND ceros_ok(9)) OR (outputA(136) AND ceros_ok(10)) OR (outputB(136) AND ceros_ok(11)) OR (outputC(136) AND ceros_ok(12)) OR (outputD(136) AND ceros_ok(13)) OR (outputE(136) AND ceros_ok(14)) OR (outputF(136) AND ceros_ok(15));
			registro_final(169) <= (output0(137) AND ceros_ok(0)) OR (output1(137) AND ceros_ok(1)) OR (output2(137) AND ceros_ok(2)) OR (output3(137) AND ceros_ok(3)) OR (output4(137) AND ceros_ok(4)) OR (output5(137) AND ceros_ok(5)) OR (output6(137) AND ceros_ok(6)) OR (output7(137) AND ceros_ok(7))OR (output8(137) AND ceros_ok(8))OR (output9(137) AND ceros_ok(9)) OR (outputA(137) AND ceros_ok(10)) OR (outputB(137) AND ceros_ok(11)) OR (outputC(137) AND ceros_ok(12)) OR (outputD(137) AND ceros_ok(13)) OR (outputE(137) AND ceros_ok(14)) OR (outputF(137) AND ceros_ok(15));
			registro_final(170) <= (output0(138) AND ceros_ok(0)) OR (output1(138) AND ceros_ok(1)) OR (output2(138) AND ceros_ok(2)) OR (output3(138) AND ceros_ok(3)) OR (output4(138) AND ceros_ok(4)) OR (output5(138) AND ceros_ok(5)) OR (output6(138) AND ceros_ok(6)) OR (output7(138) AND ceros_ok(7))OR (output8(138) AND ceros_ok(8))OR (output9(138) AND ceros_ok(9)) OR (outputA(138) AND ceros_ok(10)) OR (outputB(138) AND ceros_ok(11)) OR (outputC(138) AND ceros_ok(12)) OR (outputD(138) AND ceros_ok(13)) OR (outputE(138) AND ceros_ok(14)) OR (outputF(138) AND ceros_ok(15));
			registro_final(171) <= (output0(139) AND ceros_ok(0)) OR (output1(139) AND ceros_ok(1)) OR (output2(139) AND ceros_ok(2)) OR (output3(139) AND ceros_ok(3)) OR (output4(139) AND ceros_ok(4)) OR (output5(139) AND ceros_ok(5)) OR (output6(139) AND ceros_ok(6)) OR (output7(139) AND ceros_ok(7))OR (output8(139) AND ceros_ok(8))OR (output9(139) AND ceros_ok(9)) OR (outputA(139) AND ceros_ok(10)) OR (outputB(139) AND ceros_ok(11)) OR (outputC(139) AND ceros_ok(12)) OR (outputD(139) AND ceros_ok(13)) OR (outputE(139) AND ceros_ok(14)) OR (outputF(139) AND ceros_ok(15));
			registro_final(172) <= (output0(140) AND ceros_ok(0)) OR (output1(140) AND ceros_ok(1)) OR (output2(140) AND ceros_ok(2)) OR (output3(140) AND ceros_ok(3)) OR (output4(140) AND ceros_ok(4)) OR (output5(140) AND ceros_ok(5)) OR (output6(140) AND ceros_ok(6)) OR (output7(140) AND ceros_ok(7))OR (output8(140) AND ceros_ok(8))OR (output9(140) AND ceros_ok(9)) OR (outputA(140) AND ceros_ok(10)) OR (outputB(140) AND ceros_ok(11)) OR (outputC(140) AND ceros_ok(12)) OR (outputD(140) AND ceros_ok(13)) OR (outputE(140) AND ceros_ok(14)) OR (outputF(140) AND ceros_ok(15));
			registro_final(173) <= (output0(141) AND ceros_ok(0)) OR (output1(141) AND ceros_ok(1)) OR (output2(141) AND ceros_ok(2)) OR (output3(141) AND ceros_ok(3)) OR (output4(141) AND ceros_ok(4)) OR (output5(141) AND ceros_ok(5)) OR (output6(141) AND ceros_ok(6)) OR (output7(141) AND ceros_ok(7))OR (output8(141) AND ceros_ok(8))OR (output9(141) AND ceros_ok(9)) OR (outputA(141) AND ceros_ok(10)) OR (outputB(141) AND ceros_ok(11)) OR (outputC(141) AND ceros_ok(12)) OR (outputD(141) AND ceros_ok(13)) OR (outputE(141) AND ceros_ok(14)) OR (outputF(141) AND ceros_ok(15));
			registro_final(174) <= (output0(142) AND ceros_ok(0)) OR (output1(142) AND ceros_ok(1)) OR (output2(142) AND ceros_ok(2)) OR (output3(142) AND ceros_ok(3)) OR (output4(142) AND ceros_ok(4)) OR (output5(142) AND ceros_ok(5)) OR (output6(142) AND ceros_ok(6)) OR (output7(142) AND ceros_ok(7))OR (output8(142) AND ceros_ok(8))OR (output9(142) AND ceros_ok(9)) OR (outputA(142) AND ceros_ok(10)) OR (outputB(142) AND ceros_ok(11)) OR (outputC(142) AND ceros_ok(12)) OR (outputD(142) AND ceros_ok(13)) OR (outputE(142) AND ceros_ok(14)) OR (outputF(142) AND ceros_ok(15));
			registro_final(175) <= (output0(143) AND ceros_ok(0)) OR (output1(143) AND ceros_ok(1)) OR (output2(143) AND ceros_ok(2)) OR (output3(143) AND ceros_ok(3)) OR (output4(143) AND ceros_ok(4)) OR (output5(143) AND ceros_ok(5)) OR (output6(143) AND ceros_ok(6)) OR (output7(143) AND ceros_ok(7))OR (output8(143) AND ceros_ok(8))OR (output9(143) AND ceros_ok(9)) OR (outputA(143) AND ceros_ok(10)) OR (outputB(143) AND ceros_ok(11)) OR (outputC(143) AND ceros_ok(12)) OR (outputD(143) AND ceros_ok(13)) OR (outputE(143) AND ceros_ok(14)) OR (outputF(143) AND ceros_ok(15));
			registro_final(176) <= (output0(144) AND ceros_ok(0)) OR (output1(144) AND ceros_ok(1)) OR (output2(144) AND ceros_ok(2)) OR (output3(144) AND ceros_ok(3)) OR (output4(144) AND ceros_ok(4)) OR (output5(144) AND ceros_ok(5)) OR (output6(144) AND ceros_ok(6)) OR (output7(144) AND ceros_ok(7))OR (output8(144) AND ceros_ok(8))OR (output9(144) AND ceros_ok(9)) OR (outputA(144) AND ceros_ok(10)) OR (outputB(144) AND ceros_ok(11)) OR (outputC(144) AND ceros_ok(12)) OR (outputD(144) AND ceros_ok(13)) OR (outputE(144) AND ceros_ok(14)) OR (outputF(144) AND ceros_ok(15));
			registro_final(177) <= (output0(145) AND ceros_ok(0)) OR (output1(145) AND ceros_ok(1)) OR (output2(145) AND ceros_ok(2)) OR (output3(145) AND ceros_ok(3)) OR (output4(145) AND ceros_ok(4)) OR (output5(145) AND ceros_ok(5)) OR (output6(145) AND ceros_ok(6)) OR (output7(145) AND ceros_ok(7))OR (output8(145) AND ceros_ok(8))OR (output9(145) AND ceros_ok(9)) OR (outputA(145) AND ceros_ok(10)) OR (outputB(145) AND ceros_ok(11)) OR (outputC(145) AND ceros_ok(12)) OR (outputD(145) AND ceros_ok(13)) OR (outputE(145) AND ceros_ok(14)) OR (outputF(145) AND ceros_ok(15));
			registro_final(178) <= (output0(146) AND ceros_ok(0)) OR (output1(146) AND ceros_ok(1)) OR (output2(146) AND ceros_ok(2)) OR (output3(146) AND ceros_ok(3)) OR (output4(146) AND ceros_ok(4)) OR (output5(146) AND ceros_ok(5)) OR (output6(146) AND ceros_ok(6)) OR (output7(146) AND ceros_ok(7))OR (output8(146) AND ceros_ok(8))OR (output9(146) AND ceros_ok(9)) OR (outputA(146) AND ceros_ok(10)) OR (outputB(146) AND ceros_ok(11)) OR (outputC(146) AND ceros_ok(12)) OR (outputD(146) AND ceros_ok(13)) OR (outputE(146) AND ceros_ok(14)) OR (outputF(146) AND ceros_ok(15));
			registro_final(179) <= (output0(147) AND ceros_ok(0)) OR (output1(147) AND ceros_ok(1)) OR (output2(147) AND ceros_ok(2)) OR (output3(147) AND ceros_ok(3)) OR (output4(147) AND ceros_ok(4)) OR (output5(147) AND ceros_ok(5)) OR (output6(147) AND ceros_ok(6)) OR (output7(147) AND ceros_ok(7))OR (output8(147) AND ceros_ok(8))OR (output9(147) AND ceros_ok(9)) OR (outputA(147) AND ceros_ok(10)) OR (outputB(147) AND ceros_ok(11)) OR (outputC(147) AND ceros_ok(12)) OR (outputD(147) AND ceros_ok(13)) OR (outputE(147) AND ceros_ok(14)) OR (outputF(147) AND ceros_ok(15));
			registro_final(180) <= (output0(148) AND ceros_ok(0)) OR (output1(148) AND ceros_ok(1)) OR (output2(148) AND ceros_ok(2)) OR (output3(148) AND ceros_ok(3)) OR (output4(148) AND ceros_ok(4)) OR (output5(148) AND ceros_ok(5)) OR (output6(148) AND ceros_ok(6)) OR (output7(148) AND ceros_ok(7))OR (output8(148) AND ceros_ok(8))OR (output9(148) AND ceros_ok(9)) OR (outputA(148) AND ceros_ok(10)) OR (outputB(148) AND ceros_ok(11)) OR (outputC(148) AND ceros_ok(12)) OR (outputD(148) AND ceros_ok(13)) OR (outputE(148) AND ceros_ok(14)) OR (outputF(148) AND ceros_ok(15));
			registro_final(181) <= (output0(149) AND ceros_ok(0)) OR (output1(149) AND ceros_ok(1)) OR (output2(149) AND ceros_ok(2)) OR (output3(149) AND ceros_ok(3)) OR (output4(149) AND ceros_ok(4)) OR (output5(149) AND ceros_ok(5)) OR (output6(149) AND ceros_ok(6)) OR (output7(149) AND ceros_ok(7))OR (output8(149) AND ceros_ok(8))OR (output9(149) AND ceros_ok(9)) OR (outputA(149) AND ceros_ok(10)) OR (outputB(149) AND ceros_ok(11)) OR (outputC(149) AND ceros_ok(12)) OR (outputD(149) AND ceros_ok(13)) OR (outputE(149) AND ceros_ok(14)) OR (outputF(149) AND ceros_ok(15));
			registro_final(182) <= (output0(150) AND ceros_ok(0)) OR (output1(150) AND ceros_ok(1)) OR (output2(150) AND ceros_ok(2)) OR (output3(150) AND ceros_ok(3)) OR (output4(150) AND ceros_ok(4)) OR (output5(150) AND ceros_ok(5)) OR (output6(150) AND ceros_ok(6)) OR (output7(150) AND ceros_ok(7))OR (output8(150) AND ceros_ok(8))OR (output9(150) AND ceros_ok(9)) OR (outputA(150) AND ceros_ok(10)) OR (outputB(150) AND ceros_ok(11)) OR (outputC(150) AND ceros_ok(12)) OR (outputD(150) AND ceros_ok(13)) OR (outputE(150) AND ceros_ok(14)) OR (outputF(150) AND ceros_ok(15));
			registro_final(183) <= (output0(151) AND ceros_ok(0)) OR (output1(151) AND ceros_ok(1)) OR (output2(151) AND ceros_ok(2)) OR (output3(151) AND ceros_ok(3)) OR (output4(151) AND ceros_ok(4)) OR (output5(151) AND ceros_ok(5)) OR (output6(151) AND ceros_ok(6)) OR (output7(151) AND ceros_ok(7))OR (output8(151) AND ceros_ok(8))OR (output9(151) AND ceros_ok(9)) OR (outputA(151) AND ceros_ok(10)) OR (outputB(151) AND ceros_ok(11)) OR (outputC(151) AND ceros_ok(12)) OR (outputD(151) AND ceros_ok(13)) OR (outputE(151) AND ceros_ok(14)) OR (outputF(151) AND ceros_ok(15));
			registro_final(184) <= (output0(152) AND ceros_ok(0)) OR (output1(152) AND ceros_ok(1)) OR (output2(152) AND ceros_ok(2)) OR (output3(152) AND ceros_ok(3)) OR (output4(152) AND ceros_ok(4)) OR (output5(152) AND ceros_ok(5)) OR (output6(152) AND ceros_ok(6)) OR (output7(152) AND ceros_ok(7))OR (output8(152) AND ceros_ok(8))OR (output9(152) AND ceros_ok(9)) OR (outputA(152) AND ceros_ok(10)) OR (outputB(152) AND ceros_ok(11)) OR (outputC(152) AND ceros_ok(12)) OR (outputD(152) AND ceros_ok(13)) OR (outputE(152) AND ceros_ok(14)) OR (outputF(152) AND ceros_ok(15));
			registro_final(185) <= (output0(153) AND ceros_ok(0)) OR (output1(153) AND ceros_ok(1)) OR (output2(153) AND ceros_ok(2)) OR (output3(153) AND ceros_ok(3)) OR (output4(153) AND ceros_ok(4)) OR (output5(153) AND ceros_ok(5)) OR (output6(153) AND ceros_ok(6)) OR (output7(153) AND ceros_ok(7))OR (output8(153) AND ceros_ok(8))OR (output9(153) AND ceros_ok(9)) OR (outputA(153) AND ceros_ok(10)) OR (outputB(153) AND ceros_ok(11)) OR (outputC(153) AND ceros_ok(12)) OR (outputD(153) AND ceros_ok(13)) OR (outputE(153) AND ceros_ok(14)) OR (outputF(153) AND ceros_ok(15));
			registro_final(186) <= (output0(154) AND ceros_ok(0)) OR (output1(154) AND ceros_ok(1)) OR (output2(154) AND ceros_ok(2)) OR (output3(154) AND ceros_ok(3)) OR (output4(154) AND ceros_ok(4)) OR (output5(154) AND ceros_ok(5)) OR (output6(154) AND ceros_ok(6)) OR (output7(154) AND ceros_ok(7))OR (output8(154) AND ceros_ok(8))OR (output9(154) AND ceros_ok(9)) OR (outputA(154) AND ceros_ok(10)) OR (outputB(154) AND ceros_ok(11)) OR (outputC(154) AND ceros_ok(12)) OR (outputD(154) AND ceros_ok(13)) OR (outputE(154) AND ceros_ok(14)) OR (outputF(154) AND ceros_ok(15));
			registro_final(187) <= (output0(155) AND ceros_ok(0)) OR (output1(155) AND ceros_ok(1)) OR (output2(155) AND ceros_ok(2)) OR (output3(155) AND ceros_ok(3)) OR (output4(155) AND ceros_ok(4)) OR (output5(155) AND ceros_ok(5)) OR (output6(155) AND ceros_ok(6)) OR (output7(155) AND ceros_ok(7))OR (output8(155) AND ceros_ok(8))OR (output9(155) AND ceros_ok(9)) OR (outputA(155) AND ceros_ok(10)) OR (outputB(155) AND ceros_ok(11)) OR (outputC(155) AND ceros_ok(12)) OR (outputD(155) AND ceros_ok(13)) OR (outputE(155) AND ceros_ok(14)) OR (outputF(155) AND ceros_ok(15));
			registro_final(188) <= (output0(156) AND ceros_ok(0)) OR (output1(156) AND ceros_ok(1)) OR (output2(156) AND ceros_ok(2)) OR (output3(156) AND ceros_ok(3)) OR (output4(156) AND ceros_ok(4)) OR (output5(156) AND ceros_ok(5)) OR (output6(156) AND ceros_ok(6)) OR (output7(156) AND ceros_ok(7))OR (output8(156) AND ceros_ok(8))OR (output9(156) AND ceros_ok(9)) OR (outputA(156) AND ceros_ok(10)) OR (outputB(156) AND ceros_ok(11)) OR (outputC(156) AND ceros_ok(12)) OR (outputD(156) AND ceros_ok(13)) OR (outputE(156) AND ceros_ok(14)) OR (outputF(156) AND ceros_ok(15));
			registro_final(189) <= (output0(157) AND ceros_ok(0)) OR (output1(157) AND ceros_ok(1)) OR (output2(157) AND ceros_ok(2)) OR (output3(157) AND ceros_ok(3)) OR (output4(157) AND ceros_ok(4)) OR (output5(157) AND ceros_ok(5)) OR (output6(157) AND ceros_ok(6)) OR (output7(157) AND ceros_ok(7))OR (output8(157) AND ceros_ok(8))OR (output9(157) AND ceros_ok(9)) OR (outputA(157) AND ceros_ok(10)) OR (outputB(157) AND ceros_ok(11)) OR (outputC(157) AND ceros_ok(12)) OR (outputD(157) AND ceros_ok(13)) OR (outputE(157) AND ceros_ok(14)) OR (outputF(157) AND ceros_ok(15));
			registro_final(190) <= (output0(158) AND ceros_ok(0)) OR (output1(158) AND ceros_ok(1)) OR (output2(158) AND ceros_ok(2)) OR (output3(158) AND ceros_ok(3)) OR (output4(158) AND ceros_ok(4)) OR (output5(158) AND ceros_ok(5)) OR (output6(158) AND ceros_ok(6)) OR (output7(158) AND ceros_ok(7))OR (output8(158) AND ceros_ok(8))OR (output9(158) AND ceros_ok(9)) OR (outputA(158) AND ceros_ok(10)) OR (outputB(158) AND ceros_ok(11)) OR (outputC(158) AND ceros_ok(12)) OR (outputD(158) AND ceros_ok(13)) OR (outputE(158) AND ceros_ok(14)) OR (outputF(158) AND ceros_ok(15));
			registro_final(191) <= (output0(159) AND ceros_ok(0)) OR (output1(159) AND ceros_ok(1)) OR (output2(159) AND ceros_ok(2)) OR (output3(159) AND ceros_ok(3)) OR (output4(159) AND ceros_ok(4)) OR (output5(159) AND ceros_ok(5)) OR (output6(159) AND ceros_ok(6)) OR (output7(159) AND ceros_ok(7))OR (output8(159) AND ceros_ok(8))OR (output9(159) AND ceros_ok(9)) OR (outputA(159) AND ceros_ok(10)) OR (outputB(159) AND ceros_ok(11)) OR (outputC(159) AND ceros_ok(12)) OR (outputD(159) AND ceros_ok(13)) OR (outputE(159) AND ceros_ok(14)) OR (outputF(159) AND ceros_ok(15));
			registro_final(192) <= (output0(160) AND ceros_ok(0)) OR (output1(160) AND ceros_ok(1)) OR (output2(160) AND ceros_ok(2)) OR (output3(160) AND ceros_ok(3)) OR (output4(160) AND ceros_ok(4)) OR (output5(160) AND ceros_ok(5)) OR (output6(160) AND ceros_ok(6)) OR (output7(160) AND ceros_ok(7))OR (output8(160) AND ceros_ok(8))OR (output9(160) AND ceros_ok(9)) OR (outputA(160) AND ceros_ok(10)) OR (outputB(160) AND ceros_ok(11)) OR (outputC(160) AND ceros_ok(12)) OR (outputD(160) AND ceros_ok(13)) OR (outputE(160) AND ceros_ok(14)) OR (outputF(160) AND ceros_ok(15));
			registro_final(193) <= (output0(161) AND ceros_ok(0)) OR (output1(161) AND ceros_ok(1)) OR (output2(161) AND ceros_ok(2)) OR (output3(161) AND ceros_ok(3)) OR (output4(161) AND ceros_ok(4)) OR (output5(161) AND ceros_ok(5)) OR (output6(161) AND ceros_ok(6)) OR (output7(161) AND ceros_ok(7))OR (output8(161) AND ceros_ok(8))OR (output9(161) AND ceros_ok(9)) OR (outputA(161) AND ceros_ok(10)) OR (outputB(161) AND ceros_ok(11)) OR (outputC(161) AND ceros_ok(12)) OR (outputD(161) AND ceros_ok(13)) OR (outputE(161) AND ceros_ok(14)) OR (outputF(161) AND ceros_ok(15));
			registro_final(194) <= (output0(162) AND ceros_ok(0)) OR (output1(162) AND ceros_ok(1)) OR (output2(162) AND ceros_ok(2)) OR (output3(162) AND ceros_ok(3)) OR (output4(162) AND ceros_ok(4)) OR (output5(162) AND ceros_ok(5)) OR (output6(162) AND ceros_ok(6)) OR (output7(162) AND ceros_ok(7))OR (output8(162) AND ceros_ok(8))OR (output9(162) AND ceros_ok(9)) OR (outputA(162) AND ceros_ok(10)) OR (outputB(162) AND ceros_ok(11)) OR (outputC(162) AND ceros_ok(12)) OR (outputD(162) AND ceros_ok(13)) OR (outputE(162) AND ceros_ok(14)) OR (outputF(162) AND ceros_ok(15));
			registro_final(195) <= (output0(163) AND ceros_ok(0)) OR (output1(163) AND ceros_ok(1)) OR (output2(163) AND ceros_ok(2)) OR (output3(163) AND ceros_ok(3)) OR (output4(163) AND ceros_ok(4)) OR (output5(163) AND ceros_ok(5)) OR (output6(163) AND ceros_ok(6)) OR (output7(163) AND ceros_ok(7))OR (output8(163) AND ceros_ok(8))OR (output9(163) AND ceros_ok(9)) OR (outputA(163) AND ceros_ok(10)) OR (outputB(163) AND ceros_ok(11)) OR (outputC(163) AND ceros_ok(12)) OR (outputD(163) AND ceros_ok(13)) OR (outputE(163) AND ceros_ok(14)) OR (outputF(163) AND ceros_ok(15));
			registro_final(196) <= (output0(164) AND ceros_ok(0)) OR (output1(164) AND ceros_ok(1)) OR (output2(164) AND ceros_ok(2)) OR (output3(164) AND ceros_ok(3)) OR (output4(164) AND ceros_ok(4)) OR (output5(164) AND ceros_ok(5)) OR (output6(164) AND ceros_ok(6)) OR (output7(164) AND ceros_ok(7))OR (output8(164) AND ceros_ok(8))OR (output9(164) AND ceros_ok(9)) OR (outputA(164) AND ceros_ok(10)) OR (outputB(164) AND ceros_ok(11)) OR (outputC(164) AND ceros_ok(12)) OR (outputD(164) AND ceros_ok(13)) OR (outputE(164) AND ceros_ok(14)) OR (outputF(164) AND ceros_ok(15));
			registro_final(197) <= (output0(165) AND ceros_ok(0)) OR (output1(165) AND ceros_ok(1)) OR (output2(165) AND ceros_ok(2)) OR (output3(165) AND ceros_ok(3)) OR (output4(165) AND ceros_ok(4)) OR (output5(165) AND ceros_ok(5)) OR (output6(165) AND ceros_ok(6)) OR (output7(165) AND ceros_ok(7))OR (output8(165) AND ceros_ok(8))OR (output9(165) AND ceros_ok(9)) OR (outputA(165) AND ceros_ok(10)) OR (outputB(165) AND ceros_ok(11)) OR (outputC(165) AND ceros_ok(12)) OR (outputD(165) AND ceros_ok(13)) OR (outputE(165) AND ceros_ok(14)) OR (outputF(165) AND ceros_ok(15));
			registro_final(198) <= (output0(166) AND ceros_ok(0)) OR (output1(166) AND ceros_ok(1)) OR (output2(166) AND ceros_ok(2)) OR (output3(166) AND ceros_ok(3)) OR (output4(166) AND ceros_ok(4)) OR (output5(166) AND ceros_ok(5)) OR (output6(166) AND ceros_ok(6)) OR (output7(166) AND ceros_ok(7))OR (output8(166) AND ceros_ok(8))OR (output9(166) AND ceros_ok(9)) OR (outputA(166) AND ceros_ok(10)) OR (outputB(166) AND ceros_ok(11)) OR (outputC(166) AND ceros_ok(12)) OR (outputD(166) AND ceros_ok(13)) OR (outputE(166) AND ceros_ok(14)) OR (outputF(166) AND ceros_ok(15));
			registro_final(199) <= (output0(167) AND ceros_ok(0)) OR (output1(167) AND ceros_ok(1)) OR (output2(167) AND ceros_ok(2)) OR (output3(167) AND ceros_ok(3)) OR (output4(167) AND ceros_ok(4)) OR (output5(167) AND ceros_ok(5)) OR (output6(167) AND ceros_ok(6)) OR (output7(167) AND ceros_ok(7))OR (output8(167) AND ceros_ok(8))OR (output9(167) AND ceros_ok(9)) OR (outputA(167) AND ceros_ok(10)) OR (outputB(167) AND ceros_ok(11)) OR (outputC(167) AND ceros_ok(12)) OR (outputD(167) AND ceros_ok(13)) OR (outputE(167) AND ceros_ok(14)) OR (outputF(167) AND ceros_ok(15));
			registro_final(200) <= (output0(168) AND ceros_ok(0)) OR (output1(168) AND ceros_ok(1)) OR (output2(168) AND ceros_ok(2)) OR (output3(168) AND ceros_ok(3)) OR (output4(168) AND ceros_ok(4)) OR (output5(168) AND ceros_ok(5)) OR (output6(168) AND ceros_ok(6)) OR (output7(168) AND ceros_ok(7))OR (output8(168) AND ceros_ok(8))OR (output9(168) AND ceros_ok(9)) OR (outputA(168) AND ceros_ok(10)) OR (outputB(168) AND ceros_ok(11)) OR (outputC(168) AND ceros_ok(12)) OR (outputD(168) AND ceros_ok(13)) OR (outputE(168) AND ceros_ok(14)) OR (outputF(168) AND ceros_ok(15));
			registro_final(201) <= (output0(169) AND ceros_ok(0)) OR (output1(169) AND ceros_ok(1)) OR (output2(169) AND ceros_ok(2)) OR (output3(169) AND ceros_ok(3)) OR (output4(169) AND ceros_ok(4)) OR (output5(169) AND ceros_ok(5)) OR (output6(169) AND ceros_ok(6)) OR (output7(169) AND ceros_ok(7))OR (output8(169) AND ceros_ok(8))OR (output9(169) AND ceros_ok(9)) OR (outputA(169) AND ceros_ok(10)) OR (outputB(169) AND ceros_ok(11)) OR (outputC(169) AND ceros_ok(12)) OR (outputD(169) AND ceros_ok(13)) OR (outputE(169) AND ceros_ok(14)) OR (outputF(169) AND ceros_ok(15));
			registro_final(202) <= (output0(170) AND ceros_ok(0)) OR (output1(170) AND ceros_ok(1)) OR (output2(170) AND ceros_ok(2)) OR (output3(170) AND ceros_ok(3)) OR (output4(170) AND ceros_ok(4)) OR (output5(170) AND ceros_ok(5)) OR (output6(170) AND ceros_ok(6)) OR (output7(170) AND ceros_ok(7))OR (output8(170) AND ceros_ok(8))OR (output9(170) AND ceros_ok(9)) OR (outputA(170) AND ceros_ok(10)) OR (outputB(170) AND ceros_ok(11)) OR (outputC(170) AND ceros_ok(12)) OR (outputD(170) AND ceros_ok(13)) OR (outputE(170) AND ceros_ok(14)) OR (outputF(170) AND ceros_ok(15));
			registro_final(203) <= (output0(171) AND ceros_ok(0)) OR (output1(171) AND ceros_ok(1)) OR (output2(171) AND ceros_ok(2)) OR (output3(171) AND ceros_ok(3)) OR (output4(171) AND ceros_ok(4)) OR (output5(171) AND ceros_ok(5)) OR (output6(171) AND ceros_ok(6)) OR (output7(171) AND ceros_ok(7))OR (output8(171) AND ceros_ok(8))OR (output9(171) AND ceros_ok(9)) OR (outputA(171) AND ceros_ok(10)) OR (outputB(171) AND ceros_ok(11)) OR (outputC(171) AND ceros_ok(12)) OR (outputD(171) AND ceros_ok(13)) OR (outputE(171) AND ceros_ok(14)) OR (outputF(171) AND ceros_ok(15));
			registro_final(204) <= (output0(172) AND ceros_ok(0)) OR (output1(172) AND ceros_ok(1)) OR (output2(172) AND ceros_ok(2)) OR (output3(172) AND ceros_ok(3)) OR (output4(172) AND ceros_ok(4)) OR (output5(172) AND ceros_ok(5)) OR (output6(172) AND ceros_ok(6)) OR (output7(172) AND ceros_ok(7))OR (output8(172) AND ceros_ok(8))OR (output9(172) AND ceros_ok(9)) OR (outputA(172) AND ceros_ok(10)) OR (outputB(172) AND ceros_ok(11)) OR (outputC(172) AND ceros_ok(12)) OR (outputD(172) AND ceros_ok(13)) OR (outputE(172) AND ceros_ok(14)) OR (outputF(172) AND ceros_ok(15));
			registro_final(205) <= (output0(173) AND ceros_ok(0)) OR (output1(173) AND ceros_ok(1)) OR (output2(173) AND ceros_ok(2)) OR (output3(173) AND ceros_ok(3)) OR (output4(173) AND ceros_ok(4)) OR (output5(173) AND ceros_ok(5)) OR (output6(173) AND ceros_ok(6)) OR (output7(173) AND ceros_ok(7))OR (output8(173) AND ceros_ok(8))OR (output9(173) AND ceros_ok(9)) OR (outputA(173) AND ceros_ok(10)) OR (outputB(173) AND ceros_ok(11)) OR (outputC(173) AND ceros_ok(12)) OR (outputD(173) AND ceros_ok(13)) OR (outputE(173) AND ceros_ok(14)) OR (outputF(173) AND ceros_ok(15));
			registro_final(206) <= (output0(174) AND ceros_ok(0)) OR (output1(174) AND ceros_ok(1)) OR (output2(174) AND ceros_ok(2)) OR (output3(174) AND ceros_ok(3)) OR (output4(174) AND ceros_ok(4)) OR (output5(174) AND ceros_ok(5)) OR (output6(174) AND ceros_ok(6)) OR (output7(174) AND ceros_ok(7))OR (output8(174) AND ceros_ok(8))OR (output9(174) AND ceros_ok(9)) OR (outputA(174) AND ceros_ok(10)) OR (outputB(174) AND ceros_ok(11)) OR (outputC(174) AND ceros_ok(12)) OR (outputD(174) AND ceros_ok(13)) OR (outputE(174) AND ceros_ok(14)) OR (outputF(174) AND ceros_ok(15));
			registro_final(207) <= (output0(175) AND ceros_ok(0)) OR (output1(175) AND ceros_ok(1)) OR (output2(175) AND ceros_ok(2)) OR (output3(175) AND ceros_ok(3)) OR (output4(175) AND ceros_ok(4)) OR (output5(175) AND ceros_ok(5)) OR (output6(175) AND ceros_ok(6)) OR (output7(175) AND ceros_ok(7))OR (output8(175) AND ceros_ok(8))OR (output9(175) AND ceros_ok(9)) OR (outputA(175) AND ceros_ok(10)) OR (outputB(175) AND ceros_ok(11)) OR (outputC(175) AND ceros_ok(12)) OR (outputD(175) AND ceros_ok(13)) OR (outputE(175) AND ceros_ok(14)) OR (outputF(175) AND ceros_ok(15));
			registro_final(208) <= (output0(176) AND ceros_ok(0)) OR (output1(176) AND ceros_ok(1)) OR (output2(176) AND ceros_ok(2)) OR (output3(176) AND ceros_ok(3)) OR (output4(176) AND ceros_ok(4)) OR (output5(176) AND ceros_ok(5)) OR (output6(176) AND ceros_ok(6)) OR (output7(176) AND ceros_ok(7))OR (output8(176) AND ceros_ok(8))OR (output9(176) AND ceros_ok(9)) OR (outputA(176) AND ceros_ok(10)) OR (outputB(176) AND ceros_ok(11)) OR (outputC(176) AND ceros_ok(12)) OR (outputD(176) AND ceros_ok(13)) OR (outputE(176) AND ceros_ok(14)) OR (outputF(176) AND ceros_ok(15));
			registro_final(209) <= (output0(177) AND ceros_ok(0)) OR (output1(177) AND ceros_ok(1)) OR (output2(177) AND ceros_ok(2)) OR (output3(177) AND ceros_ok(3)) OR (output4(177) AND ceros_ok(4)) OR (output5(177) AND ceros_ok(5)) OR (output6(177) AND ceros_ok(6)) OR (output7(177) AND ceros_ok(7))OR (output8(177) AND ceros_ok(8))OR (output9(177) AND ceros_ok(9)) OR (outputA(177) AND ceros_ok(10)) OR (outputB(177) AND ceros_ok(11)) OR (outputC(177) AND ceros_ok(12)) OR (outputD(177) AND ceros_ok(13)) OR (outputE(177) AND ceros_ok(14)) OR (outputF(177) AND ceros_ok(15));
			registro_final(210) <= (output0(178) AND ceros_ok(0)) OR (output1(178) AND ceros_ok(1)) OR (output2(178) AND ceros_ok(2)) OR (output3(178) AND ceros_ok(3)) OR (output4(178) AND ceros_ok(4)) OR (output5(178) AND ceros_ok(5)) OR (output6(178) AND ceros_ok(6)) OR (output7(178) AND ceros_ok(7))OR (output8(178) AND ceros_ok(8))OR (output9(178) AND ceros_ok(9)) OR (outputA(178) AND ceros_ok(10)) OR (outputB(178) AND ceros_ok(11)) OR (outputC(178) AND ceros_ok(12)) OR (outputD(178) AND ceros_ok(13)) OR (outputE(178) AND ceros_ok(14)) OR (outputF(178) AND ceros_ok(15));
			registro_final(211) <= (output0(179) AND ceros_ok(0)) OR (output1(179) AND ceros_ok(1)) OR (output2(179) AND ceros_ok(2)) OR (output3(179) AND ceros_ok(3)) OR (output4(179) AND ceros_ok(4)) OR (output5(179) AND ceros_ok(5)) OR (output6(179) AND ceros_ok(6)) OR (output7(179) AND ceros_ok(7))OR (output8(179) AND ceros_ok(8))OR (output9(179) AND ceros_ok(9)) OR (outputA(179) AND ceros_ok(10)) OR (outputB(179) AND ceros_ok(11)) OR (outputC(179) AND ceros_ok(12)) OR (outputD(179) AND ceros_ok(13)) OR (outputE(179) AND ceros_ok(14)) OR (outputF(179) AND ceros_ok(15));
			registro_final(212) <= (output0(180) AND ceros_ok(0)) OR (output1(180) AND ceros_ok(1)) OR (output2(180) AND ceros_ok(2)) OR (output3(180) AND ceros_ok(3)) OR (output4(180) AND ceros_ok(4)) OR (output5(180) AND ceros_ok(5)) OR (output6(180) AND ceros_ok(6)) OR (output7(180) AND ceros_ok(7))OR (output8(180) AND ceros_ok(8))OR (output9(180) AND ceros_ok(9)) OR (outputA(180) AND ceros_ok(10)) OR (outputB(180) AND ceros_ok(11)) OR (outputC(180) AND ceros_ok(12)) OR (outputD(180) AND ceros_ok(13)) OR (outputE(180) AND ceros_ok(14)) OR (outputF(180) AND ceros_ok(15));
			registro_final(213) <= (output0(181) AND ceros_ok(0)) OR (output1(181) AND ceros_ok(1)) OR (output2(181) AND ceros_ok(2)) OR (output3(181) AND ceros_ok(3)) OR (output4(181) AND ceros_ok(4)) OR (output5(181) AND ceros_ok(5)) OR (output6(181) AND ceros_ok(6)) OR (output7(181) AND ceros_ok(7))OR (output8(181) AND ceros_ok(8))OR (output9(181) AND ceros_ok(9)) OR (outputA(181) AND ceros_ok(10)) OR (outputB(181) AND ceros_ok(11)) OR (outputC(181) AND ceros_ok(12)) OR (outputD(181) AND ceros_ok(13)) OR (outputE(181) AND ceros_ok(14)) OR (outputF(181) AND ceros_ok(15));
			registro_final(214) <= (output0(182) AND ceros_ok(0)) OR (output1(182) AND ceros_ok(1)) OR (output2(182) AND ceros_ok(2)) OR (output3(182) AND ceros_ok(3)) OR (output4(182) AND ceros_ok(4)) OR (output5(182) AND ceros_ok(5)) OR (output6(182) AND ceros_ok(6)) OR (output7(182) AND ceros_ok(7))OR (output8(182) AND ceros_ok(8))OR (output9(182) AND ceros_ok(9)) OR (outputA(182) AND ceros_ok(10)) OR (outputB(182) AND ceros_ok(11)) OR (outputC(182) AND ceros_ok(12)) OR (outputD(182) AND ceros_ok(13)) OR (outputE(182) AND ceros_ok(14)) OR (outputF(182) AND ceros_ok(15));
			registro_final(215) <= (output0(183) AND ceros_ok(0)) OR (output1(183) AND ceros_ok(1)) OR (output2(183) AND ceros_ok(2)) OR (output3(183) AND ceros_ok(3)) OR (output4(183) AND ceros_ok(4)) OR (output5(183) AND ceros_ok(5)) OR (output6(183) AND ceros_ok(6)) OR (output7(183) AND ceros_ok(7))OR (output8(183) AND ceros_ok(8))OR (output9(183) AND ceros_ok(9)) OR (outputA(183) AND ceros_ok(10)) OR (outputB(183) AND ceros_ok(11)) OR (outputC(183) AND ceros_ok(12)) OR (outputD(183) AND ceros_ok(13)) OR (outputE(183) AND ceros_ok(14)) OR (outputF(183) AND ceros_ok(15));
			registro_final(216) <= (output0(184) AND ceros_ok(0)) OR (output1(184) AND ceros_ok(1)) OR (output2(184) AND ceros_ok(2)) OR (output3(184) AND ceros_ok(3)) OR (output4(184) AND ceros_ok(4)) OR (output5(184) AND ceros_ok(5)) OR (output6(184) AND ceros_ok(6)) OR (output7(184) AND ceros_ok(7))OR (output8(184) AND ceros_ok(8))OR (output9(184) AND ceros_ok(9)) OR (outputA(184) AND ceros_ok(10)) OR (outputB(184) AND ceros_ok(11)) OR (outputC(184) AND ceros_ok(12)) OR (outputD(184) AND ceros_ok(13)) OR (outputE(184) AND ceros_ok(14)) OR (outputF(184) AND ceros_ok(15));
			registro_final(217) <= (output0(185) AND ceros_ok(0)) OR (output1(185) AND ceros_ok(1)) OR (output2(185) AND ceros_ok(2)) OR (output3(185) AND ceros_ok(3)) OR (output4(185) AND ceros_ok(4)) OR (output5(185) AND ceros_ok(5)) OR (output6(185) AND ceros_ok(6)) OR (output7(185) AND ceros_ok(7))OR (output8(185) AND ceros_ok(8))OR (output9(185) AND ceros_ok(9)) OR (outputA(185) AND ceros_ok(10)) OR (outputB(185) AND ceros_ok(11)) OR (outputC(185) AND ceros_ok(12)) OR (outputD(185) AND ceros_ok(13)) OR (outputE(185) AND ceros_ok(14)) OR (outputF(185) AND ceros_ok(15));
			registro_final(218) <= (output0(186) AND ceros_ok(0)) OR (output1(186) AND ceros_ok(1)) OR (output2(186) AND ceros_ok(2)) OR (output3(186) AND ceros_ok(3)) OR (output4(186) AND ceros_ok(4)) OR (output5(186) AND ceros_ok(5)) OR (output6(186) AND ceros_ok(6)) OR (output7(186) AND ceros_ok(7))OR (output8(186) AND ceros_ok(8))OR (output9(186) AND ceros_ok(9)) OR (outputA(186) AND ceros_ok(10)) OR (outputB(186) AND ceros_ok(11)) OR (outputC(186) AND ceros_ok(12)) OR (outputD(186) AND ceros_ok(13)) OR (outputE(186) AND ceros_ok(14)) OR (outputF(186) AND ceros_ok(15));
			registro_final(219) <= (output0(187) AND ceros_ok(0)) OR (output1(187) AND ceros_ok(1)) OR (output2(187) AND ceros_ok(2)) OR (output3(187) AND ceros_ok(3)) OR (output4(187) AND ceros_ok(4)) OR (output5(187) AND ceros_ok(5)) OR (output6(187) AND ceros_ok(6)) OR (output7(187) AND ceros_ok(7))OR (output8(187) AND ceros_ok(8))OR (output9(187) AND ceros_ok(9)) OR (outputA(187) AND ceros_ok(10)) OR (outputB(187) AND ceros_ok(11)) OR (outputC(187) AND ceros_ok(12)) OR (outputD(187) AND ceros_ok(13)) OR (outputE(187) AND ceros_ok(14)) OR (outputF(187) AND ceros_ok(15));
			registro_final(220) <= (output0(188) AND ceros_ok(0)) OR (output1(188) AND ceros_ok(1)) OR (output2(188) AND ceros_ok(2)) OR (output3(188) AND ceros_ok(3)) OR (output4(188) AND ceros_ok(4)) OR (output5(188) AND ceros_ok(5)) OR (output6(188) AND ceros_ok(6)) OR (output7(188) AND ceros_ok(7))OR (output8(188) AND ceros_ok(8))OR (output9(188) AND ceros_ok(9)) OR (outputA(188) AND ceros_ok(10)) OR (outputB(188) AND ceros_ok(11)) OR (outputC(188) AND ceros_ok(12)) OR (outputD(188) AND ceros_ok(13)) OR (outputE(188) AND ceros_ok(14)) OR (outputF(188) AND ceros_ok(15));
			registro_final(221) <= (output0(189) AND ceros_ok(0)) OR (output1(189) AND ceros_ok(1)) OR (output2(189) AND ceros_ok(2)) OR (output3(189) AND ceros_ok(3)) OR (output4(189) AND ceros_ok(4)) OR (output5(189) AND ceros_ok(5)) OR (output6(189) AND ceros_ok(6)) OR (output7(189) AND ceros_ok(7))OR (output8(189) AND ceros_ok(8))OR (output9(189) AND ceros_ok(9)) OR (outputA(189) AND ceros_ok(10)) OR (outputB(189) AND ceros_ok(11)) OR (outputC(189) AND ceros_ok(12)) OR (outputD(189) AND ceros_ok(13)) OR (outputE(189) AND ceros_ok(14)) OR (outputF(189) AND ceros_ok(15));
			registro_final(222) <= (output0(190) AND ceros_ok(0)) OR (output1(190) AND ceros_ok(1)) OR (output2(190) AND ceros_ok(2)) OR (output3(190) AND ceros_ok(3)) OR (output4(190) AND ceros_ok(4)) OR (output5(190) AND ceros_ok(5)) OR (output6(190) AND ceros_ok(6)) OR (output7(190) AND ceros_ok(7))OR (output8(190) AND ceros_ok(8))OR (output9(190) AND ceros_ok(9)) OR (outputA(190) AND ceros_ok(10)) OR (outputB(190) AND ceros_ok(11)) OR (outputC(190) AND ceros_ok(12)) OR (outputD(190) AND ceros_ok(13)) OR (outputE(190) AND ceros_ok(14)) OR (outputF(190) AND ceros_ok(15));
			registro_final(223) <= (output0(191) AND ceros_ok(0)) OR (output1(191) AND ceros_ok(1)) OR (output2(191) AND ceros_ok(2)) OR (output3(191) AND ceros_ok(3)) OR (output4(191) AND ceros_ok(4)) OR (output5(191) AND ceros_ok(5)) OR (output6(191) AND ceros_ok(6)) OR (output7(191) AND ceros_ok(7))OR (output8(191) AND ceros_ok(8))OR (output9(191) AND ceros_ok(9)) OR (outputA(191) AND ceros_ok(10)) OR (outputB(191) AND ceros_ok(11)) OR (outputC(191) AND ceros_ok(12)) OR (outputD(191) AND ceros_ok(13)) OR (outputE(191) AND ceros_ok(14)) OR (outputF(191) AND ceros_ok(15));
			registro_final(224) <= (output0(192) AND ceros_ok(0)) OR (output1(192) AND ceros_ok(1)) OR (output2(192) AND ceros_ok(2)) OR (output3(192) AND ceros_ok(3)) OR (output4(192) AND ceros_ok(4)) OR (output5(192) AND ceros_ok(5)) OR (output6(192) AND ceros_ok(6)) OR (output7(192) AND ceros_ok(7))OR (output8(192) AND ceros_ok(8))OR (output9(192) AND ceros_ok(9)) OR (outputA(192) AND ceros_ok(10)) OR (outputB(192) AND ceros_ok(11)) OR (outputC(192) AND ceros_ok(12)) OR (outputD(192) AND ceros_ok(13)) OR (outputE(192) AND ceros_ok(14)) OR (outputF(192) AND ceros_ok(15));
			registro_final(225) <= (output0(193) AND ceros_ok(0)) OR (output1(193) AND ceros_ok(1)) OR (output2(193) AND ceros_ok(2)) OR (output3(193) AND ceros_ok(3)) OR (output4(193) AND ceros_ok(4)) OR (output5(193) AND ceros_ok(5)) OR (output6(193) AND ceros_ok(6)) OR (output7(193) AND ceros_ok(7))OR (output8(193) AND ceros_ok(8))OR (output9(193) AND ceros_ok(9)) OR (outputA(193) AND ceros_ok(10)) OR (outputB(193) AND ceros_ok(11)) OR (outputC(193) AND ceros_ok(12)) OR (outputD(193) AND ceros_ok(13)) OR (outputE(193) AND ceros_ok(14)) OR (outputF(193) AND ceros_ok(15));
			registro_final(226) <= (output0(194) AND ceros_ok(0)) OR (output1(194) AND ceros_ok(1)) OR (output2(194) AND ceros_ok(2)) OR (output3(194) AND ceros_ok(3)) OR (output4(194) AND ceros_ok(4)) OR (output5(194) AND ceros_ok(5)) OR (output6(194) AND ceros_ok(6)) OR (output7(194) AND ceros_ok(7))OR (output8(194) AND ceros_ok(8))OR (output9(194) AND ceros_ok(9)) OR (outputA(194) AND ceros_ok(10)) OR (outputB(194) AND ceros_ok(11)) OR (outputC(194) AND ceros_ok(12)) OR (outputD(194) AND ceros_ok(13)) OR (outputE(194) AND ceros_ok(14)) OR (outputF(194) AND ceros_ok(15));
			registro_final(227) <= (output0(195) AND ceros_ok(0)) OR (output1(195) AND ceros_ok(1)) OR (output2(195) AND ceros_ok(2)) OR (output3(195) AND ceros_ok(3)) OR (output4(195) AND ceros_ok(4)) OR (output5(195) AND ceros_ok(5)) OR (output6(195) AND ceros_ok(6)) OR (output7(195) AND ceros_ok(7))OR (output8(195) AND ceros_ok(8))OR (output9(195) AND ceros_ok(9)) OR (outputA(195) AND ceros_ok(10)) OR (outputB(195) AND ceros_ok(11)) OR (outputC(195) AND ceros_ok(12)) OR (outputD(195) AND ceros_ok(13)) OR (outputE(195) AND ceros_ok(14)) OR (outputF(195) AND ceros_ok(15));
			registro_final(228) <= (output0(196) AND ceros_ok(0)) OR (output1(196) AND ceros_ok(1)) OR (output2(196) AND ceros_ok(2)) OR (output3(196) AND ceros_ok(3)) OR (output4(196) AND ceros_ok(4)) OR (output5(196) AND ceros_ok(5)) OR (output6(196) AND ceros_ok(6)) OR (output7(196) AND ceros_ok(7))OR (output8(196) AND ceros_ok(8))OR (output9(196) AND ceros_ok(9)) OR (outputA(196) AND ceros_ok(10)) OR (outputB(196) AND ceros_ok(11)) OR (outputC(196) AND ceros_ok(12)) OR (outputD(196) AND ceros_ok(13)) OR (outputE(196) AND ceros_ok(14)) OR (outputF(196) AND ceros_ok(15));
			registro_final(229) <= (output0(197) AND ceros_ok(0)) OR (output1(197) AND ceros_ok(1)) OR (output2(197) AND ceros_ok(2)) OR (output3(197) AND ceros_ok(3)) OR (output4(197) AND ceros_ok(4)) OR (output5(197) AND ceros_ok(5)) OR (output6(197) AND ceros_ok(6)) OR (output7(197) AND ceros_ok(7))OR (output8(197) AND ceros_ok(8))OR (output9(197) AND ceros_ok(9)) OR (outputA(197) AND ceros_ok(10)) OR (outputB(197) AND ceros_ok(11)) OR (outputC(197) AND ceros_ok(12)) OR (outputD(197) AND ceros_ok(13)) OR (outputE(197) AND ceros_ok(14)) OR (outputF(197) AND ceros_ok(15));
			registro_final(230) <= (output0(198) AND ceros_ok(0)) OR (output1(198) AND ceros_ok(1)) OR (output2(198) AND ceros_ok(2)) OR (output3(198) AND ceros_ok(3)) OR (output4(198) AND ceros_ok(4)) OR (output5(198) AND ceros_ok(5)) OR (output6(198) AND ceros_ok(6)) OR (output7(198) AND ceros_ok(7))OR (output8(198) AND ceros_ok(8))OR (output9(198) AND ceros_ok(9)) OR (outputA(198) AND ceros_ok(10)) OR (outputB(198) AND ceros_ok(11)) OR (outputC(198) AND ceros_ok(12)) OR (outputD(198) AND ceros_ok(13)) OR (outputE(198) AND ceros_ok(14)) OR (outputF(198) AND ceros_ok(15));
			registro_final(231) <= (output0(199) AND ceros_ok(0)) OR (output1(199) AND ceros_ok(1)) OR (output2(199) AND ceros_ok(2)) OR (output3(199) AND ceros_ok(3)) OR (output4(199) AND ceros_ok(4)) OR (output5(199) AND ceros_ok(5)) OR (output6(199) AND ceros_ok(6)) OR (output7(199) AND ceros_ok(7))OR (output8(199) AND ceros_ok(8))OR (output9(199) AND ceros_ok(9)) OR (outputA(199) AND ceros_ok(10)) OR (outputB(199) AND ceros_ok(11)) OR (outputC(199) AND ceros_ok(12)) OR (outputD(199) AND ceros_ok(13)) OR (outputE(199) AND ceros_ok(14)) OR (outputF(199) AND ceros_ok(15));
			registro_final(232) <= (output0(200) AND ceros_ok(0)) OR (output1(200) AND ceros_ok(1)) OR (output2(200) AND ceros_ok(2)) OR (output3(200) AND ceros_ok(3)) OR (output4(200) AND ceros_ok(4)) OR (output5(200) AND ceros_ok(5)) OR (output6(200) AND ceros_ok(6)) OR (output7(200) AND ceros_ok(7))OR (output8(200) AND ceros_ok(8))OR (output9(200) AND ceros_ok(9)) OR (outputA(200) AND ceros_ok(10)) OR (outputB(200) AND ceros_ok(11)) OR (outputC(200) AND ceros_ok(12)) OR (outputD(200) AND ceros_ok(13)) OR (outputE(200) AND ceros_ok(14)) OR (outputF(200) AND ceros_ok(15));
			registro_final(233) <= (output0(201) AND ceros_ok(0)) OR (output1(201) AND ceros_ok(1)) OR (output2(201) AND ceros_ok(2)) OR (output3(201) AND ceros_ok(3)) OR (output4(201) AND ceros_ok(4)) OR (output5(201) AND ceros_ok(5)) OR (output6(201) AND ceros_ok(6)) OR (output7(201) AND ceros_ok(7))OR (output8(201) AND ceros_ok(8))OR (output9(201) AND ceros_ok(9)) OR (outputA(201) AND ceros_ok(10)) OR (outputB(201) AND ceros_ok(11)) OR (outputC(201) AND ceros_ok(12)) OR (outputD(201) AND ceros_ok(13)) OR (outputE(201) AND ceros_ok(14)) OR (outputF(201) AND ceros_ok(15));
			registro_final(234) <= (output0(202) AND ceros_ok(0)) OR (output1(202) AND ceros_ok(1)) OR (output2(202) AND ceros_ok(2)) OR (output3(202) AND ceros_ok(3)) OR (output4(202) AND ceros_ok(4)) OR (output5(202) AND ceros_ok(5)) OR (output6(202) AND ceros_ok(6)) OR (output7(202) AND ceros_ok(7))OR (output8(202) AND ceros_ok(8))OR (output9(202) AND ceros_ok(9)) OR (outputA(202) AND ceros_ok(10)) OR (outputB(202) AND ceros_ok(11)) OR (outputC(202) AND ceros_ok(12)) OR (outputD(202) AND ceros_ok(13)) OR (outputE(202) AND ceros_ok(14)) OR (outputF(202) AND ceros_ok(15));
			registro_final(235) <= (output0(203) AND ceros_ok(0)) OR (output1(203) AND ceros_ok(1)) OR (output2(203) AND ceros_ok(2)) OR (output3(203) AND ceros_ok(3)) OR (output4(203) AND ceros_ok(4)) OR (output5(203) AND ceros_ok(5)) OR (output6(203) AND ceros_ok(6)) OR (output7(203) AND ceros_ok(7))OR (output8(203) AND ceros_ok(8))OR (output9(203) AND ceros_ok(9)) OR (outputA(203) AND ceros_ok(10)) OR (outputB(203) AND ceros_ok(11)) OR (outputC(203) AND ceros_ok(12)) OR (outputD(203) AND ceros_ok(13)) OR (outputE(203) AND ceros_ok(14)) OR (outputF(203) AND ceros_ok(15));
			registro_final(236) <= (output0(204) AND ceros_ok(0)) OR (output1(204) AND ceros_ok(1)) OR (output2(204) AND ceros_ok(2)) OR (output3(204) AND ceros_ok(3)) OR (output4(204) AND ceros_ok(4)) OR (output5(204) AND ceros_ok(5)) OR (output6(204) AND ceros_ok(6)) OR (output7(204) AND ceros_ok(7))OR (output8(204) AND ceros_ok(8))OR (output9(204) AND ceros_ok(9)) OR (outputA(204) AND ceros_ok(10)) OR (outputB(204) AND ceros_ok(11)) OR (outputC(204) AND ceros_ok(12)) OR (outputD(204) AND ceros_ok(13)) OR (outputE(204) AND ceros_ok(14)) OR (outputF(204) AND ceros_ok(15));
			registro_final(237) <= (output0(205) AND ceros_ok(0)) OR (output1(205) AND ceros_ok(1)) OR (output2(205) AND ceros_ok(2)) OR (output3(205) AND ceros_ok(3)) OR (output4(205) AND ceros_ok(4)) OR (output5(205) AND ceros_ok(5)) OR (output6(205) AND ceros_ok(6)) OR (output7(205) AND ceros_ok(7))OR (output8(205) AND ceros_ok(8))OR (output9(205) AND ceros_ok(9)) OR (outputA(205) AND ceros_ok(10)) OR (outputB(205) AND ceros_ok(11)) OR (outputC(205) AND ceros_ok(12)) OR (outputD(205) AND ceros_ok(13)) OR (outputE(205) AND ceros_ok(14)) OR (outputF(205) AND ceros_ok(15));
			registro_final(238) <= (output0(206) AND ceros_ok(0)) OR (output1(206) AND ceros_ok(1)) OR (output2(206) AND ceros_ok(2)) OR (output3(206) AND ceros_ok(3)) OR (output4(206) AND ceros_ok(4)) OR (output5(206) AND ceros_ok(5)) OR (output6(206) AND ceros_ok(6)) OR (output7(206) AND ceros_ok(7))OR (output8(206) AND ceros_ok(8))OR (output9(206) AND ceros_ok(9)) OR (outputA(206) AND ceros_ok(10)) OR (outputB(206) AND ceros_ok(11)) OR (outputC(206) AND ceros_ok(12)) OR (outputD(206) AND ceros_ok(13)) OR (outputE(206) AND ceros_ok(14)) OR (outputF(206) AND ceros_ok(15));
			registro_final(239) <= (output0(207) AND ceros_ok(0)) OR (output1(207) AND ceros_ok(1)) OR (output2(207) AND ceros_ok(2)) OR (output3(207) AND ceros_ok(3)) OR (output4(207) AND ceros_ok(4)) OR (output5(207) AND ceros_ok(5)) OR (output6(207) AND ceros_ok(6)) OR (output7(207) AND ceros_ok(7))OR (output8(207) AND ceros_ok(8))OR (output9(207) AND ceros_ok(9)) OR (outputA(207) AND ceros_ok(10)) OR (outputB(207) AND ceros_ok(11)) OR (outputC(207) AND ceros_ok(12)) OR (outputD(207) AND ceros_ok(13)) OR (outputE(207) AND ceros_ok(14)) OR (outputF(207) AND ceros_ok(15));
			registro_final(240) <= (output0(208) AND ceros_ok(0)) OR (output1(208) AND ceros_ok(1)) OR (output2(208) AND ceros_ok(2)) OR (output3(208) AND ceros_ok(3)) OR (output4(208) AND ceros_ok(4)) OR (output5(208) AND ceros_ok(5)) OR (output6(208) AND ceros_ok(6)) OR (output7(208) AND ceros_ok(7))OR (output8(208) AND ceros_ok(8))OR (output9(208) AND ceros_ok(9)) OR (outputA(208) AND ceros_ok(10)) OR (outputB(208) AND ceros_ok(11)) OR (outputC(208) AND ceros_ok(12)) OR (outputD(208) AND ceros_ok(13)) OR (outputE(208) AND ceros_ok(14)) OR (outputF(208) AND ceros_ok(15));
			registro_final(241) <= (output0(209) AND ceros_ok(0)) OR (output1(209) AND ceros_ok(1)) OR (output2(209) AND ceros_ok(2)) OR (output3(209) AND ceros_ok(3)) OR (output4(209) AND ceros_ok(4)) OR (output5(209) AND ceros_ok(5)) OR (output6(209) AND ceros_ok(6)) OR (output7(209) AND ceros_ok(7))OR (output8(209) AND ceros_ok(8))OR (output9(209) AND ceros_ok(9)) OR (outputA(209) AND ceros_ok(10)) OR (outputB(209) AND ceros_ok(11)) OR (outputC(209) AND ceros_ok(12)) OR (outputD(209) AND ceros_ok(13)) OR (outputE(209) AND ceros_ok(14)) OR (outputF(209) AND ceros_ok(15));
			registro_final(242) <= (output0(210) AND ceros_ok(0)) OR (output1(210) AND ceros_ok(1)) OR (output2(210) AND ceros_ok(2)) OR (output3(210) AND ceros_ok(3)) OR (output4(210) AND ceros_ok(4)) OR (output5(210) AND ceros_ok(5)) OR (output6(210) AND ceros_ok(6)) OR (output7(210) AND ceros_ok(7))OR (output8(210) AND ceros_ok(8))OR (output9(210) AND ceros_ok(9)) OR (outputA(210) AND ceros_ok(10)) OR (outputB(210) AND ceros_ok(11)) OR (outputC(210) AND ceros_ok(12)) OR (outputD(210) AND ceros_ok(13)) OR (outputE(210) AND ceros_ok(14)) OR (outputF(210) AND ceros_ok(15));
			registro_final(243) <= (output0(211) AND ceros_ok(0)) OR (output1(211) AND ceros_ok(1)) OR (output2(211) AND ceros_ok(2)) OR (output3(211) AND ceros_ok(3)) OR (output4(211) AND ceros_ok(4)) OR (output5(211) AND ceros_ok(5)) OR (output6(211) AND ceros_ok(6)) OR (output7(211) AND ceros_ok(7))OR (output8(211) AND ceros_ok(8))OR (output9(211) AND ceros_ok(9)) OR (outputA(211) AND ceros_ok(10)) OR (outputB(211) AND ceros_ok(11)) OR (outputC(211) AND ceros_ok(12)) OR (outputD(211) AND ceros_ok(13)) OR (outputE(211) AND ceros_ok(14)) OR (outputF(211) AND ceros_ok(15));
			registro_final(244) <= (output0(212) AND ceros_ok(0)) OR (output1(212) AND ceros_ok(1)) OR (output2(212) AND ceros_ok(2)) OR (output3(212) AND ceros_ok(3)) OR (output4(212) AND ceros_ok(4)) OR (output5(212) AND ceros_ok(5)) OR (output6(212) AND ceros_ok(6)) OR (output7(212) AND ceros_ok(7))OR (output8(212) AND ceros_ok(8))OR (output9(212) AND ceros_ok(9)) OR (outputA(212) AND ceros_ok(10)) OR (outputB(212) AND ceros_ok(11)) OR (outputC(212) AND ceros_ok(12)) OR (outputD(212) AND ceros_ok(13)) OR (outputE(212) AND ceros_ok(14)) OR (outputF(212) AND ceros_ok(15));
			registro_final(245) <= (output0(213) AND ceros_ok(0)) OR (output1(213) AND ceros_ok(1)) OR (output2(213) AND ceros_ok(2)) OR (output3(213) AND ceros_ok(3)) OR (output4(213) AND ceros_ok(4)) OR (output5(213) AND ceros_ok(5)) OR (output6(213) AND ceros_ok(6)) OR (output7(213) AND ceros_ok(7))OR (output8(213) AND ceros_ok(8))OR (output9(213) AND ceros_ok(9)) OR (outputA(213) AND ceros_ok(10)) OR (outputB(213) AND ceros_ok(11)) OR (outputC(213) AND ceros_ok(12)) OR (outputD(213) AND ceros_ok(13)) OR (outputE(213) AND ceros_ok(14)) OR (outputF(213) AND ceros_ok(15));
			registro_final(246) <= (output0(214) AND ceros_ok(0)) OR (output1(214) AND ceros_ok(1)) OR (output2(214) AND ceros_ok(2)) OR (output3(214) AND ceros_ok(3)) OR (output4(214) AND ceros_ok(4)) OR (output5(214) AND ceros_ok(5)) OR (output6(214) AND ceros_ok(6)) OR (output7(214) AND ceros_ok(7))OR (output8(214) AND ceros_ok(8))OR (output9(214) AND ceros_ok(9)) OR (outputA(214) AND ceros_ok(10)) OR (outputB(214) AND ceros_ok(11)) OR (outputC(214) AND ceros_ok(12)) OR (outputD(214) AND ceros_ok(13)) OR (outputE(214) AND ceros_ok(14)) OR (outputF(214) AND ceros_ok(15));
			registro_final(247) <= (output0(215) AND ceros_ok(0)) OR (output1(215) AND ceros_ok(1)) OR (output2(215) AND ceros_ok(2)) OR (output3(215) AND ceros_ok(3)) OR (output4(215) AND ceros_ok(4)) OR (output5(215) AND ceros_ok(5)) OR (output6(215) AND ceros_ok(6)) OR (output7(215) AND ceros_ok(7))OR (output8(215) AND ceros_ok(8))OR (output9(215) AND ceros_ok(9)) OR (outputA(215) AND ceros_ok(10)) OR (outputB(215) AND ceros_ok(11)) OR (outputC(215) AND ceros_ok(12)) OR (outputD(215) AND ceros_ok(13)) OR (outputE(215) AND ceros_ok(14)) OR (outputF(215) AND ceros_ok(15));
			registro_final(248) <= (output0(216) AND ceros_ok(0)) OR (output1(216) AND ceros_ok(1)) OR (output2(216) AND ceros_ok(2)) OR (output3(216) AND ceros_ok(3)) OR (output4(216) AND ceros_ok(4)) OR (output5(216) AND ceros_ok(5)) OR (output6(216) AND ceros_ok(6)) OR (output7(216) AND ceros_ok(7))OR (output8(216) AND ceros_ok(8))OR (output9(216) AND ceros_ok(9)) OR (outputA(216) AND ceros_ok(10)) OR (outputB(216) AND ceros_ok(11)) OR (outputC(216) AND ceros_ok(12)) OR (outputD(216) AND ceros_ok(13)) OR (outputE(216) AND ceros_ok(14)) OR (outputF(216) AND ceros_ok(15));
			registro_final(249) <= (output0(217) AND ceros_ok(0)) OR (output1(217) AND ceros_ok(1)) OR (output2(217) AND ceros_ok(2)) OR (output3(217) AND ceros_ok(3)) OR (output4(217) AND ceros_ok(4)) OR (output5(217) AND ceros_ok(5)) OR (output6(217) AND ceros_ok(6)) OR (output7(217) AND ceros_ok(7))OR (output8(217) AND ceros_ok(8))OR (output9(217) AND ceros_ok(9)) OR (outputA(217) AND ceros_ok(10)) OR (outputB(217) AND ceros_ok(11)) OR (outputC(217) AND ceros_ok(12)) OR (outputD(217) AND ceros_ok(13)) OR (outputE(217) AND ceros_ok(14)) OR (outputF(217) AND ceros_ok(15));
			registro_final(250) <= (output0(218) AND ceros_ok(0)) OR (output1(218) AND ceros_ok(1)) OR (output2(218) AND ceros_ok(2)) OR (output3(218) AND ceros_ok(3)) OR (output4(218) AND ceros_ok(4)) OR (output5(218) AND ceros_ok(5)) OR (output6(218) AND ceros_ok(6)) OR (output7(218) AND ceros_ok(7))OR (output8(218) AND ceros_ok(8))OR (output9(218) AND ceros_ok(9)) OR (outputA(218) AND ceros_ok(10)) OR (outputB(218) AND ceros_ok(11)) OR (outputC(218) AND ceros_ok(12)) OR (outputD(218) AND ceros_ok(13)) OR (outputE(218) AND ceros_ok(14)) OR (outputF(218) AND ceros_ok(15));
			registro_final(251) <= (output0(219) AND ceros_ok(0)) OR (output1(219) AND ceros_ok(1)) OR (output2(219) AND ceros_ok(2)) OR (output3(219) AND ceros_ok(3)) OR (output4(219) AND ceros_ok(4)) OR (output5(219) AND ceros_ok(5)) OR (output6(219) AND ceros_ok(6)) OR (output7(219) AND ceros_ok(7))OR (output8(219) AND ceros_ok(8))OR (output9(219) AND ceros_ok(9)) OR (outputA(219) AND ceros_ok(10)) OR (outputB(219) AND ceros_ok(11)) OR (outputC(219) AND ceros_ok(12)) OR (outputD(219) AND ceros_ok(13)) OR (outputE(219) AND ceros_ok(14)) OR (outputF(219) AND ceros_ok(15));
			registro_final(252) <= (output0(220) AND ceros_ok(0)) OR (output1(220) AND ceros_ok(1)) OR (output2(220) AND ceros_ok(2)) OR (output3(220) AND ceros_ok(3)) OR (output4(220) AND ceros_ok(4)) OR (output5(220) AND ceros_ok(5)) OR (output6(220) AND ceros_ok(6)) OR (output7(220) AND ceros_ok(7))OR (output8(220) AND ceros_ok(8))OR (output9(220) AND ceros_ok(9)) OR (outputA(220) AND ceros_ok(10)) OR (outputB(220) AND ceros_ok(11)) OR (outputC(220) AND ceros_ok(12)) OR (outputD(220) AND ceros_ok(13)) OR (outputE(220) AND ceros_ok(14)) OR (outputF(220) AND ceros_ok(15));
			registro_final(253) <= (output0(221) AND ceros_ok(0)) OR (output1(221) AND ceros_ok(1)) OR (output2(221) AND ceros_ok(2)) OR (output3(221) AND ceros_ok(3)) OR (output4(221) AND ceros_ok(4)) OR (output5(221) AND ceros_ok(5)) OR (output6(221) AND ceros_ok(6)) OR (output7(221) AND ceros_ok(7))OR (output8(221) AND ceros_ok(8))OR (output9(221) AND ceros_ok(9)) OR (outputA(221) AND ceros_ok(10)) OR (outputB(221) AND ceros_ok(11)) OR (outputC(221) AND ceros_ok(12)) OR (outputD(221) AND ceros_ok(13)) OR (outputE(221) AND ceros_ok(14)) OR (outputF(221) AND ceros_ok(15));
			registro_final(254) <= (output0(222) AND ceros_ok(0)) OR (output1(222) AND ceros_ok(1)) OR (output2(222) AND ceros_ok(2)) OR (output3(222) AND ceros_ok(3)) OR (output4(222) AND ceros_ok(4)) OR (output5(222) AND ceros_ok(5)) OR (output6(222) AND ceros_ok(6)) OR (output7(222) AND ceros_ok(7))OR (output8(222) AND ceros_ok(8))OR (output9(222) AND ceros_ok(9)) OR (outputA(222) AND ceros_ok(10)) OR (outputB(222) AND ceros_ok(11)) OR (outputC(222) AND ceros_ok(12)) OR (outputD(222) AND ceros_ok(13)) OR (outputE(222) AND ceros_ok(14)) OR (outputF(222) AND ceros_ok(15));
			registro_final(255) <= (output0(223) AND ceros_ok(0)) OR (output1(223) AND ceros_ok(1)) OR (output2(223) AND ceros_ok(2)) OR (output3(223) AND ceros_ok(3)) OR (output4(223) AND ceros_ok(4)) OR (output5(223) AND ceros_ok(5)) OR (output6(223) AND ceros_ok(6)) OR (output7(223) AND ceros_ok(7))OR (output8(223) AND ceros_ok(8))OR (output9(223) AND ceros_ok(9)) OR (outputA(223) AND ceros_ok(10)) OR (outputB(223) AND ceros_ok(11)) OR (outputC(223) AND ceros_ok(12)) OR (outputD(223) AND ceros_ok(13)) OR (outputE(223) AND ceros_ok(14)) OR (outputF(223) AND ceros_ok(15));
			registro_final(256) <= (output0(224) AND ceros_ok(0)) OR (output1(224) AND ceros_ok(1)) OR (output2(224) AND ceros_ok(2)) OR (output3(224) AND ceros_ok(3)) OR (output4(224) AND ceros_ok(4)) OR (output5(224) AND ceros_ok(5)) OR (output6(224) AND ceros_ok(6)) OR (output7(224) AND ceros_ok(7))OR (output8(224) AND ceros_ok(8))OR (output9(224) AND ceros_ok(9)) OR (outputA(224) AND ceros_ok(10)) OR (outputB(224) AND ceros_ok(11)) OR (outputC(224) AND ceros_ok(12)) OR (outputD(224) AND ceros_ok(13)) OR (outputE(224) AND ceros_ok(14)) OR (outputF(224) AND ceros_ok(15));
			registro_final(257) <= (output0(225) AND ceros_ok(0)) OR (output1(225) AND ceros_ok(1)) OR (output2(225) AND ceros_ok(2)) OR (output3(225) AND ceros_ok(3)) OR (output4(225) AND ceros_ok(4)) OR (output5(225) AND ceros_ok(5)) OR (output6(225) AND ceros_ok(6)) OR (output7(225) AND ceros_ok(7))OR (output8(225) AND ceros_ok(8))OR (output9(225) AND ceros_ok(9)) OR (outputA(225) AND ceros_ok(10)) OR (outputB(225) AND ceros_ok(11)) OR (outputC(225) AND ceros_ok(12)) OR (outputD(225) AND ceros_ok(13)) OR (outputE(225) AND ceros_ok(14)) OR (outputF(225) AND ceros_ok(15));
			registro_final(258) <= (output0(226) AND ceros_ok(0)) OR (output1(226) AND ceros_ok(1)) OR (output2(226) AND ceros_ok(2)) OR (output3(226) AND ceros_ok(3)) OR (output4(226) AND ceros_ok(4)) OR (output5(226) AND ceros_ok(5)) OR (output6(226) AND ceros_ok(6)) OR (output7(226) AND ceros_ok(7))OR (output8(226) AND ceros_ok(8))OR (output9(226) AND ceros_ok(9)) OR (outputA(226) AND ceros_ok(10)) OR (outputB(226) AND ceros_ok(11)) OR (outputC(226) AND ceros_ok(12)) OR (outputD(226) AND ceros_ok(13)) OR (outputE(226) AND ceros_ok(14)) OR (outputF(226) AND ceros_ok(15));
			registro_final(259) <= (output0(227) AND ceros_ok(0)) OR (output1(227) AND ceros_ok(1)) OR (output2(227) AND ceros_ok(2)) OR (output3(227) AND ceros_ok(3)) OR (output4(227) AND ceros_ok(4)) OR (output5(227) AND ceros_ok(5)) OR (output6(227) AND ceros_ok(6)) OR (output7(227) AND ceros_ok(7))OR (output8(227) AND ceros_ok(8))OR (output9(227) AND ceros_ok(9)) OR (outputA(227) AND ceros_ok(10)) OR (outputB(227) AND ceros_ok(11)) OR (outputC(227) AND ceros_ok(12)) OR (outputD(227) AND ceros_ok(13)) OR (outputE(227) AND ceros_ok(14)) OR (outputF(227) AND ceros_ok(15));
			registro_final(260) <= (output0(228) AND ceros_ok(0)) OR (output1(228) AND ceros_ok(1)) OR (output2(228) AND ceros_ok(2)) OR (output3(228) AND ceros_ok(3)) OR (output4(228) AND ceros_ok(4)) OR (output5(228) AND ceros_ok(5)) OR (output6(228) AND ceros_ok(6)) OR (output7(228) AND ceros_ok(7))OR (output8(228) AND ceros_ok(8))OR (output9(228) AND ceros_ok(9)) OR (outputA(228) AND ceros_ok(10)) OR (outputB(228) AND ceros_ok(11)) OR (outputC(228) AND ceros_ok(12)) OR (outputD(228) AND ceros_ok(13)) OR (outputE(228) AND ceros_ok(14)) OR (outputF(228) AND ceros_ok(15));
			registro_final(261) <= (output0(229) AND ceros_ok(0)) OR (output1(229) AND ceros_ok(1)) OR (output2(229) AND ceros_ok(2)) OR (output3(229) AND ceros_ok(3)) OR (output4(229) AND ceros_ok(4)) OR (output5(229) AND ceros_ok(5)) OR (output6(229) AND ceros_ok(6)) OR (output7(229) AND ceros_ok(7))OR (output8(229) AND ceros_ok(8))OR (output9(229) AND ceros_ok(9)) OR (outputA(229) AND ceros_ok(10)) OR (outputB(229) AND ceros_ok(11)) OR (outputC(229) AND ceros_ok(12)) OR (outputD(229) AND ceros_ok(13)) OR (outputE(229) AND ceros_ok(14)) OR (outputF(229) AND ceros_ok(15));
			registro_final(262) <= (output0(230) AND ceros_ok(0)) OR (output1(230) AND ceros_ok(1)) OR (output2(230) AND ceros_ok(2)) OR (output3(230) AND ceros_ok(3)) OR (output4(230) AND ceros_ok(4)) OR (output5(230) AND ceros_ok(5)) OR (output6(230) AND ceros_ok(6)) OR (output7(230) AND ceros_ok(7))OR (output8(230) AND ceros_ok(8))OR (output9(230) AND ceros_ok(9)) OR (outputA(230) AND ceros_ok(10)) OR (outputB(230) AND ceros_ok(11)) OR (outputC(230) AND ceros_ok(12)) OR (outputD(230) AND ceros_ok(13)) OR (outputE(230) AND ceros_ok(14)) OR (outputF(230) AND ceros_ok(15));
			registro_final(263) <= (output0(231) AND ceros_ok(0)) OR (output1(231) AND ceros_ok(1)) OR (output2(231) AND ceros_ok(2)) OR (output3(231) AND ceros_ok(3)) OR (output4(231) AND ceros_ok(4)) OR (output5(231) AND ceros_ok(5)) OR (output6(231) AND ceros_ok(6)) OR (output7(231) AND ceros_ok(7))OR (output8(231) AND ceros_ok(8))OR (output9(231) AND ceros_ok(9)) OR (outputA(231) AND ceros_ok(10)) OR (outputB(231) AND ceros_ok(11)) OR (outputC(231) AND ceros_ok(12)) OR (outputD(231) AND ceros_ok(13)) OR (outputE(231) AND ceros_ok(14)) OR (outputF(231) AND ceros_ok(15));
			registro_final(264) <= (output0(232) AND ceros_ok(0)) OR (output1(232) AND ceros_ok(1)) OR (output2(232) AND ceros_ok(2)) OR (output3(232) AND ceros_ok(3)) OR (output4(232) AND ceros_ok(4)) OR (output5(232) AND ceros_ok(5)) OR (output6(232) AND ceros_ok(6)) OR (output7(232) AND ceros_ok(7))OR (output8(232) AND ceros_ok(8))OR (output9(232) AND ceros_ok(9)) OR (outputA(232) AND ceros_ok(10)) OR (outputB(232) AND ceros_ok(11)) OR (outputC(232) AND ceros_ok(12)) OR (outputD(232) AND ceros_ok(13)) OR (outputE(232) AND ceros_ok(14)) OR (outputF(232) AND ceros_ok(15));
			registro_final(265) <= (output0(233) AND ceros_ok(0)) OR (output1(233) AND ceros_ok(1)) OR (output2(233) AND ceros_ok(2)) OR (output3(233) AND ceros_ok(3)) OR (output4(233) AND ceros_ok(4)) OR (output5(233) AND ceros_ok(5)) OR (output6(233) AND ceros_ok(6)) OR (output7(233) AND ceros_ok(7))OR (output8(233) AND ceros_ok(8))OR (output9(233) AND ceros_ok(9)) OR (outputA(233) AND ceros_ok(10)) OR (outputB(233) AND ceros_ok(11)) OR (outputC(233) AND ceros_ok(12)) OR (outputD(233) AND ceros_ok(13)) OR (outputE(233) AND ceros_ok(14)) OR (outputF(233) AND ceros_ok(15));
			registro_final(266) <= (output0(234) AND ceros_ok(0)) OR (output1(234) AND ceros_ok(1)) OR (output2(234) AND ceros_ok(2)) OR (output3(234) AND ceros_ok(3)) OR (output4(234) AND ceros_ok(4)) OR (output5(234) AND ceros_ok(5)) OR (output6(234) AND ceros_ok(6)) OR (output7(234) AND ceros_ok(7))OR (output8(234) AND ceros_ok(8))OR (output9(234) AND ceros_ok(9)) OR (outputA(234) AND ceros_ok(10)) OR (outputB(234) AND ceros_ok(11)) OR (outputC(234) AND ceros_ok(12)) OR (outputD(234) AND ceros_ok(13)) OR (outputE(234) AND ceros_ok(14)) OR (outputF(234) AND ceros_ok(15));
			registro_final(267) <= (output0(235) AND ceros_ok(0)) OR (output1(235) AND ceros_ok(1)) OR (output2(235) AND ceros_ok(2)) OR (output3(235) AND ceros_ok(3)) OR (output4(235) AND ceros_ok(4)) OR (output5(235) AND ceros_ok(5)) OR (output6(235) AND ceros_ok(6)) OR (output7(235) AND ceros_ok(7))OR (output8(235) AND ceros_ok(8))OR (output9(235) AND ceros_ok(9)) OR (outputA(235) AND ceros_ok(10)) OR (outputB(235) AND ceros_ok(11)) OR (outputC(235) AND ceros_ok(12)) OR (outputD(235) AND ceros_ok(13)) OR (outputE(235) AND ceros_ok(14)) OR (outputF(235) AND ceros_ok(15));
			registro_final(268) <= (output0(236) AND ceros_ok(0)) OR (output1(236) AND ceros_ok(1)) OR (output2(236) AND ceros_ok(2)) OR (output3(236) AND ceros_ok(3)) OR (output4(236) AND ceros_ok(4)) OR (output5(236) AND ceros_ok(5)) OR (output6(236) AND ceros_ok(6)) OR (output7(236) AND ceros_ok(7))OR (output8(236) AND ceros_ok(8))OR (output9(236) AND ceros_ok(9)) OR (outputA(236) AND ceros_ok(10)) OR (outputB(236) AND ceros_ok(11)) OR (outputC(236) AND ceros_ok(12)) OR (outputD(236) AND ceros_ok(13)) OR (outputE(236) AND ceros_ok(14)) OR (outputF(236) AND ceros_ok(15));
			registro_final(269) <= (output0(237) AND ceros_ok(0)) OR (output1(237) AND ceros_ok(1)) OR (output2(237) AND ceros_ok(2)) OR (output3(237) AND ceros_ok(3)) OR (output4(237) AND ceros_ok(4)) OR (output5(237) AND ceros_ok(5)) OR (output6(237) AND ceros_ok(6)) OR (output7(237) AND ceros_ok(7))OR (output8(237) AND ceros_ok(8))OR (output9(237) AND ceros_ok(9)) OR (outputA(237) AND ceros_ok(10)) OR (outputB(237) AND ceros_ok(11)) OR (outputC(237) AND ceros_ok(12)) OR (outputD(237) AND ceros_ok(13)) OR (outputE(237) AND ceros_ok(14)) OR (outputF(237) AND ceros_ok(15));
			registro_final(270) <= (output0(238) AND ceros_ok(0)) OR (output1(238) AND ceros_ok(1)) OR (output2(238) AND ceros_ok(2)) OR (output3(238) AND ceros_ok(3)) OR (output4(238) AND ceros_ok(4)) OR (output5(238) AND ceros_ok(5)) OR (output6(238) AND ceros_ok(6)) OR (output7(238) AND ceros_ok(7))OR (output8(238) AND ceros_ok(8))OR (output9(238) AND ceros_ok(9)) OR (outputA(238) AND ceros_ok(10)) OR (outputB(238) AND ceros_ok(11)) OR (outputC(238) AND ceros_ok(12)) OR (outputD(238) AND ceros_ok(13)) OR (outputE(238) AND ceros_ok(14)) OR (outputF(238) AND ceros_ok(15));
			registro_final(271) <= (output0(239) AND ceros_ok(0)) OR (output1(239) AND ceros_ok(1)) OR (output2(239) AND ceros_ok(2)) OR (output3(239) AND ceros_ok(3)) OR (output4(239) AND ceros_ok(4)) OR (output5(239) AND ceros_ok(5)) OR (output6(239) AND ceros_ok(6)) OR (output7(239) AND ceros_ok(7))OR (output8(239) AND ceros_ok(8))OR (output9(239) AND ceros_ok(9)) OR (outputA(239) AND ceros_ok(10)) OR (outputB(239) AND ceros_ok(11)) OR (outputC(239) AND ceros_ok(12)) OR (outputD(239) AND ceros_ok(13)) OR (outputE(239) AND ceros_ok(14)) OR (outputF(239) AND ceros_ok(15));
			registro_final(272) <= (output0(240) AND ceros_ok(0)) OR (output1(240) AND ceros_ok(1)) OR (output2(240) AND ceros_ok(2)) OR (output3(240) AND ceros_ok(3)) OR (output4(240) AND ceros_ok(4)) OR (output5(240) AND ceros_ok(5)) OR (output6(240) AND ceros_ok(6)) OR (output7(240) AND ceros_ok(7))OR (output8(240) AND ceros_ok(8))OR (output9(240) AND ceros_ok(9)) OR (outputA(240) AND ceros_ok(10)) OR (outputB(240) AND ceros_ok(11)) OR (outputC(240) AND ceros_ok(12)) OR (outputD(240) AND ceros_ok(13)) OR (outputE(240) AND ceros_ok(14)) OR (outputF(240) AND ceros_ok(15));
			registro_final(273) <= (output0(241) AND ceros_ok(0)) OR (output1(241) AND ceros_ok(1)) OR (output2(241) AND ceros_ok(2)) OR (output3(241) AND ceros_ok(3)) OR (output4(241) AND ceros_ok(4)) OR (output5(241) AND ceros_ok(5)) OR (output6(241) AND ceros_ok(6)) OR (output7(241) AND ceros_ok(7))OR (output8(241) AND ceros_ok(8))OR (output9(241) AND ceros_ok(9)) OR (outputA(241) AND ceros_ok(10)) OR (outputB(241) AND ceros_ok(11)) OR (outputC(241) AND ceros_ok(12)) OR (outputD(241) AND ceros_ok(13)) OR (outputE(241) AND ceros_ok(14)) OR (outputF(241) AND ceros_ok(15));
			registro_final(274) <= (output0(242) AND ceros_ok(0)) OR (output1(242) AND ceros_ok(1)) OR (output2(242) AND ceros_ok(2)) OR (output3(242) AND ceros_ok(3)) OR (output4(242) AND ceros_ok(4)) OR (output5(242) AND ceros_ok(5)) OR (output6(242) AND ceros_ok(6)) OR (output7(242) AND ceros_ok(7))OR (output8(242) AND ceros_ok(8))OR (output9(242) AND ceros_ok(9)) OR (outputA(242) AND ceros_ok(10)) OR (outputB(242) AND ceros_ok(11)) OR (outputC(242) AND ceros_ok(12)) OR (outputD(242) AND ceros_ok(13)) OR (outputE(242) AND ceros_ok(14)) OR (outputF(242) AND ceros_ok(15));
			registro_final(275) <= (output0(243) AND ceros_ok(0)) OR (output1(243) AND ceros_ok(1)) OR (output2(243) AND ceros_ok(2)) OR (output3(243) AND ceros_ok(3)) OR (output4(243) AND ceros_ok(4)) OR (output5(243) AND ceros_ok(5)) OR (output6(243) AND ceros_ok(6)) OR (output7(243) AND ceros_ok(7))OR (output8(243) AND ceros_ok(8))OR (output9(243) AND ceros_ok(9)) OR (outputA(243) AND ceros_ok(10)) OR (outputB(243) AND ceros_ok(11)) OR (outputC(243) AND ceros_ok(12)) OR (outputD(243) AND ceros_ok(13)) OR (outputE(243) AND ceros_ok(14)) OR (outputF(243) AND ceros_ok(15));
			registro_final(276) <= (output0(244) AND ceros_ok(0)) OR (output1(244) AND ceros_ok(1)) OR (output2(244) AND ceros_ok(2)) OR (output3(244) AND ceros_ok(3)) OR (output4(244) AND ceros_ok(4)) OR (output5(244) AND ceros_ok(5)) OR (output6(244) AND ceros_ok(6)) OR (output7(244) AND ceros_ok(7))OR (output8(244) AND ceros_ok(8))OR (output9(244) AND ceros_ok(9)) OR (outputA(244) AND ceros_ok(10)) OR (outputB(244) AND ceros_ok(11)) OR (outputC(244) AND ceros_ok(12)) OR (outputD(244) AND ceros_ok(13)) OR (outputE(244) AND ceros_ok(14)) OR (outputF(244) AND ceros_ok(15));
			registro_final(277) <= (output0(245) AND ceros_ok(0)) OR (output1(245) AND ceros_ok(1)) OR (output2(245) AND ceros_ok(2)) OR (output3(245) AND ceros_ok(3)) OR (output4(245) AND ceros_ok(4)) OR (output5(245) AND ceros_ok(5)) OR (output6(245) AND ceros_ok(6)) OR (output7(245) AND ceros_ok(7))OR (output8(245) AND ceros_ok(8))OR (output9(245) AND ceros_ok(9)) OR (outputA(245) AND ceros_ok(10)) OR (outputB(245) AND ceros_ok(11)) OR (outputC(245) AND ceros_ok(12)) OR (outputD(245) AND ceros_ok(13)) OR (outputE(245) AND ceros_ok(14)) OR (outputF(245) AND ceros_ok(15));
			registro_final(278) <= (output0(246) AND ceros_ok(0)) OR (output1(246) AND ceros_ok(1)) OR (output2(246) AND ceros_ok(2)) OR (output3(246) AND ceros_ok(3)) OR (output4(246) AND ceros_ok(4)) OR (output5(246) AND ceros_ok(5)) OR (output6(246) AND ceros_ok(6)) OR (output7(246) AND ceros_ok(7))OR (output8(246) AND ceros_ok(8))OR (output9(246) AND ceros_ok(9)) OR (outputA(246) AND ceros_ok(10)) OR (outputB(246) AND ceros_ok(11)) OR (outputC(246) AND ceros_ok(12)) OR (outputD(246) AND ceros_ok(13)) OR (outputE(246) AND ceros_ok(14)) OR (outputF(246) AND ceros_ok(15));
			registro_final(279) <= (output0(247) AND ceros_ok(0)) OR (output1(247) AND ceros_ok(1)) OR (output2(247) AND ceros_ok(2)) OR (output3(247) AND ceros_ok(3)) OR (output4(247) AND ceros_ok(4)) OR (output5(247) AND ceros_ok(5)) OR (output6(247) AND ceros_ok(6)) OR (output7(247) AND ceros_ok(7))OR (output8(247) AND ceros_ok(8))OR (output9(247) AND ceros_ok(9)) OR (outputA(247) AND ceros_ok(10)) OR (outputB(247) AND ceros_ok(11)) OR (outputC(247) AND ceros_ok(12)) OR (outputD(247) AND ceros_ok(13)) OR (outputE(247) AND ceros_ok(14)) OR (outputF(247) AND ceros_ok(15));
			registro_final(280) <= (output0(248) AND ceros_ok(0)) OR (output1(248) AND ceros_ok(1)) OR (output2(248) AND ceros_ok(2)) OR (output3(248) AND ceros_ok(3)) OR (output4(248) AND ceros_ok(4)) OR (output5(248) AND ceros_ok(5)) OR (output6(248) AND ceros_ok(6)) OR (output7(248) AND ceros_ok(7))OR (output8(248) AND ceros_ok(8))OR (output9(248) AND ceros_ok(9)) OR (outputA(248) AND ceros_ok(10)) OR (outputB(248) AND ceros_ok(11)) OR (outputC(248) AND ceros_ok(12)) OR (outputD(248) AND ceros_ok(13)) OR (outputE(248) AND ceros_ok(14)) OR (outputF(248) AND ceros_ok(15));
			registro_final(281) <= (output0(249) AND ceros_ok(0)) OR (output1(249) AND ceros_ok(1)) OR (output2(249) AND ceros_ok(2)) OR (output3(249) AND ceros_ok(3)) OR (output4(249) AND ceros_ok(4)) OR (output5(249) AND ceros_ok(5)) OR (output6(249) AND ceros_ok(6)) OR (output7(249) AND ceros_ok(7))OR (output8(249) AND ceros_ok(8))OR (output9(249) AND ceros_ok(9)) OR (outputA(249) AND ceros_ok(10)) OR (outputB(249) AND ceros_ok(11)) OR (outputC(249) AND ceros_ok(12)) OR (outputD(249) AND ceros_ok(13)) OR (outputE(249) AND ceros_ok(14)) OR (outputF(249) AND ceros_ok(15));
			registro_final(282) <= (output0(250) AND ceros_ok(0)) OR (output1(250) AND ceros_ok(1)) OR (output2(250) AND ceros_ok(2)) OR (output3(250) AND ceros_ok(3)) OR (output4(250) AND ceros_ok(4)) OR (output5(250) AND ceros_ok(5)) OR (output6(250) AND ceros_ok(6)) OR (output7(250) AND ceros_ok(7))OR (output8(250) AND ceros_ok(8))OR (output9(250) AND ceros_ok(9)) OR (outputA(250) AND ceros_ok(10)) OR (outputB(250) AND ceros_ok(11)) OR (outputC(250) AND ceros_ok(12)) OR (outputD(250) AND ceros_ok(13)) OR (outputE(250) AND ceros_ok(14)) OR (outputF(250) AND ceros_ok(15));
			registro_final(283) <= (output0(251) AND ceros_ok(0)) OR (output1(251) AND ceros_ok(1)) OR (output2(251) AND ceros_ok(2)) OR (output3(251) AND ceros_ok(3)) OR (output4(251) AND ceros_ok(4)) OR (output5(251) AND ceros_ok(5)) OR (output6(251) AND ceros_ok(6)) OR (output7(251) AND ceros_ok(7))OR (output8(251) AND ceros_ok(8))OR (output9(251) AND ceros_ok(9)) OR (outputA(251) AND ceros_ok(10)) OR (outputB(251) AND ceros_ok(11)) OR (outputC(251) AND ceros_ok(12)) OR (outputD(251) AND ceros_ok(13)) OR (outputE(251) AND ceros_ok(14)) OR (outputF(251) AND ceros_ok(15));
			registro_final(284) <= (output0(252) AND ceros_ok(0)) OR (output1(252) AND ceros_ok(1)) OR (output2(252) AND ceros_ok(2)) OR (output3(252) AND ceros_ok(3)) OR (output4(252) AND ceros_ok(4)) OR (output5(252) AND ceros_ok(5)) OR (output6(252) AND ceros_ok(6)) OR (output7(252) AND ceros_ok(7))OR (output8(252) AND ceros_ok(8))OR (output9(252) AND ceros_ok(9)) OR (outputA(252) AND ceros_ok(10)) OR (outputB(252) AND ceros_ok(11)) OR (outputC(252) AND ceros_ok(12)) OR (outputD(252) AND ceros_ok(13)) OR (outputE(252) AND ceros_ok(14)) OR (outputF(252) AND ceros_ok(15));
			registro_final(285) <= (output0(253) AND ceros_ok(0)) OR (output1(253) AND ceros_ok(1)) OR (output2(253) AND ceros_ok(2)) OR (output3(253) AND ceros_ok(3)) OR (output4(253) AND ceros_ok(4)) OR (output5(253) AND ceros_ok(5)) OR (output6(253) AND ceros_ok(6)) OR (output7(253) AND ceros_ok(7))OR (output8(253) AND ceros_ok(8))OR (output9(253) AND ceros_ok(9)) OR (outputA(253) AND ceros_ok(10)) OR (outputB(253) AND ceros_ok(11)) OR (outputC(253) AND ceros_ok(12)) OR (outputD(253) AND ceros_ok(13)) OR (outputE(253) AND ceros_ok(14)) OR (outputF(253) AND ceros_ok(15));
			registro_final(286) <= (output0(254) AND ceros_ok(0)) OR (output1(254) AND ceros_ok(1)) OR (output2(254) AND ceros_ok(2)) OR (output3(254) AND ceros_ok(3)) OR (output4(254) AND ceros_ok(4)) OR (output5(254) AND ceros_ok(5)) OR (output6(254) AND ceros_ok(6)) OR (output7(254) AND ceros_ok(7))OR (output8(254) AND ceros_ok(8))OR (output9(254) AND ceros_ok(9)) OR (outputA(254) AND ceros_ok(10)) OR (outputB(254) AND ceros_ok(11)) OR (outputC(254) AND ceros_ok(12)) OR (outputD(254) AND ceros_ok(13)) OR (outputE(254) AND ceros_ok(14)) OR (outputF(254) AND ceros_ok(15));
			registro_final(287) <= (output0(255) AND ceros_ok(0)) OR (output1(255) AND ceros_ok(1)) OR (output2(255) AND ceros_ok(2)) OR (output3(255) AND ceros_ok(3)) OR (output4(255) AND ceros_ok(4)) OR (output5(255) AND ceros_ok(5)) OR (output6(255) AND ceros_ok(6)) OR (output7(255) AND ceros_ok(7))OR (output8(255) AND ceros_ok(8))OR (output9(255) AND ceros_ok(9)) OR (outputA(255) AND ceros_ok(10)) OR (outputB(255) AND ceros_ok(11)) OR (outputC(255) AND ceros_ok(12)) OR (outputD(255) AND ceros_ok(13)) OR (outputE(255) AND ceros_ok(14)) OR (outputF(255) AND ceros_ok(15));

			END IF;
		END IF;
	END PROCESS;
END ARCHITECTURE Output_selArchh;