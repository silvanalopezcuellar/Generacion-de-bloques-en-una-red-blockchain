LIBRARY ieee;
USE ieee.STD_LOGIC_1164.all;
USE ieee.numeric_std.all;
-------------------------------------
ENTITY RAM IS
	GENERIC (Xmax : integer:= 511;
				Ymax : integer:= 16 ;
				halfL : integer);
	PORT(	 	clk		  		: IN 	STD_ULOGIC;
				wr_en		  		: IN 	STD_ULOGIC;
				data_in	  		: IN 	STD_ULOGIC;
				bloques			: IN 	INTEGER ;
				fin_mensaje		: IN 	STD_ULOGIC;
				--read
				row_rd_addr 	: IN INTEGER ;
				column_rd_addr : IN INTEGER ;
				--write
				row_wr_addr 	: IN INTEGER :=0;
				column_wr_addr : IN INTEGER :=0;
				finalByte		: OUT STD_ULOGIC_VECTOR (halfL-1 DOWNTO 0);
				data_out			: OUT STD_ULOGIC_VECTOR (511 DOWNTO 0)
		  );
END RAM;
--------------------------------------
ARCHITECTURE behavioral OF RAM IS
	TYPE data 		IS ARRAY (Ymax DOWNTO 0) OF STD_ULOGIC;
	TYPE mem_type 	IS ARRAY (Xmax DOWNTO 0) OF data;
	SIGNAL 	mem : mem_type := (others => (others => '0'));
	
BEGIN
	--write process
	write_process: PROCESS(clk)
	BEGIN
		IF (rising_edge(clk)) THEN
			IF(fin_mensaje='1' AND bloques>=1) THEN
			
				finalByte(5) <= mem(509)(bloques-1);
				finalByte(4) <= mem(508)(bloques-1);
				finalByte(3) <= mem(507)(bloques-1);
				finalByte(2) <= mem(506)(bloques-1);
				finalByte(1) <= mem(505)(bloques-1);
				finalByte(0) <= mem(504)(bloques-1);
				
			END IF;
			
		IF(wr_en = '1' AND column_wr_addr>=0 AND row_wr_addr>=0) THEN
				mem(row_wr_addr)(column_wr_addr)<= data_in;
		END IF;
		 	
								data_out(7)  <=mem(511)(column_rd_addr);
								data_out(6)  <=mem(510)(column_rd_addr);
								data_out(5)  <=mem(509)(column_rd_addr);
								data_out(4)  <=mem(508)(column_rd_addr);
								data_out(3)  <=mem(507)(column_rd_addr);
								data_out(2)  <=mem(506)(column_rd_addr);
								data_out(1)  <=mem(505)(column_rd_addr);
								data_out(0)  <=mem(504)(column_rd_addr);
								data_out(15) <=mem(503)(column_rd_addr);
								data_out(14) <=mem(502)(column_rd_addr);
								data_out(13) <=mem(501)(column_rd_addr);
								data_out(12) <=mem(500)(column_rd_addr);
								data_out(11) <=mem(499)(column_rd_addr);
								data_out(10) <=mem(498)(column_rd_addr);
								data_out(9)  <=mem(497)(column_rd_addr);
								data_out(8)  <=mem(496)(column_rd_addr);
								data_out(23) <=mem(495)(column_rd_addr);
								data_out(22) <=mem(494)(column_rd_addr);
								data_out(21) <=mem(493)(column_rd_addr);
								data_out(20) <=mem(492)(column_rd_addr);
								data_out(19) <=mem(491)(column_rd_addr);
								data_out(18) <=mem(490)(column_rd_addr);
								data_out(17) <=mem(489)(column_rd_addr);
								data_out(16) <=mem(488)(column_rd_addr);
								data_out(31) <=mem(487)(column_rd_addr);
								data_out(30) <=mem(486)(column_rd_addr);
								data_out(29) <=mem(485)(column_rd_addr);
								data_out(28) <=mem(484)(column_rd_addr);
								data_out(27) <=mem(483)(column_rd_addr);
								data_out(26) <=mem(482)(column_rd_addr);
								data_out(25) <=mem(481)(column_rd_addr);
								data_out(24) <=mem(480)(column_rd_addr);
								data_out(39) <=mem(479)(column_rd_addr);
								data_out(38) <=mem(478)(column_rd_addr);
								data_out(37) <=mem(477)(column_rd_addr);
								data_out(36) <=mem(476)(column_rd_addr);
								data_out(35) <=mem(475)(column_rd_addr);
								data_out(34) <=mem(474)(column_rd_addr);
								data_out(33) <=mem(473)(column_rd_addr);
								data_out(32) <=mem(472)(column_rd_addr);
								data_out(47) <=mem(471)(column_rd_addr);
								data_out(46) <=mem(470)(column_rd_addr);
								data_out(45) <=mem(469)(column_rd_addr);
								data_out(44) <=mem(468)(column_rd_addr);
								data_out(43) <=mem(467)(column_rd_addr);
								data_out(42) <=mem(466)(column_rd_addr);
								data_out(41) <=mem(465)(column_rd_addr);
								data_out(40) <=mem(464)(column_rd_addr);
								data_out(55) <=mem(463)(column_rd_addr);
								data_out(54) <=mem(462)(column_rd_addr);
								data_out(53) <=mem(461)(column_rd_addr);
								data_out(52) <=mem(460)(column_rd_addr);
								data_out(51) <=mem(459)(column_rd_addr);
								data_out(50) <=mem(458)(column_rd_addr);
								data_out(49) <=mem(457)(column_rd_addr);
								data_out(48) <=mem(456)(column_rd_addr);
								data_out(63) <=mem(455)(column_rd_addr);
								data_out(62) <=mem(454)(column_rd_addr);
								data_out(61) <=mem(453)(column_rd_addr);
								data_out(60) <=mem(452)(column_rd_addr);
								data_out(59) <=mem(451)(column_rd_addr);
								data_out(58) <=mem(450)(column_rd_addr);
								data_out(57) <=mem(449)(column_rd_addr);
								data_out(56) <=mem(448)(column_rd_addr);
								data_out(71) <=mem(447)(column_rd_addr);
								data_out(70) <=mem(446)(column_rd_addr);
								data_out(69) <=mem(445)(column_rd_addr);
								data_out(68) <=mem(444)(column_rd_addr);
								data_out(67) <=mem(443)(column_rd_addr);
								data_out(66) <=mem(442)(column_rd_addr);
								data_out(65) <=mem(441)(column_rd_addr);
								data_out(64) <=mem(440)(column_rd_addr);
								data_out(79) <=mem(439)(column_rd_addr);
								data_out(78) <=mem(438)(column_rd_addr);
								data_out(77) <=mem(437)(column_rd_addr);
								data_out(76) <=mem(436)(column_rd_addr);
								data_out(75) <=mem(435)(column_rd_addr);
								data_out(74) <=mem(434)(column_rd_addr);
								data_out(73) <=mem(433)(column_rd_addr);
								data_out(72) <=mem(432)(column_rd_addr);
								data_out(87) <=mem(431)(column_rd_addr);
								data_out(86) <=mem(430)(column_rd_addr);
								data_out(85) <=mem(429)(column_rd_addr);
								data_out(84) <=mem(428)(column_rd_addr);
								data_out(83) <=mem(427)(column_rd_addr);
								data_out(82) <=mem(426)(column_rd_addr);
								data_out(81) <=mem(425)(column_rd_addr);
								data_out(80) <=mem(424)(column_rd_addr);
								data_out(95) <=mem(423)(column_rd_addr);
								data_out(94) <=mem(422)(column_rd_addr);
								data_out(93) <=mem(421)(column_rd_addr);
								data_out(92) <=mem(420)(column_rd_addr);
								data_out(91) <=mem(419)(column_rd_addr);
								data_out(90) <=mem(418)(column_rd_addr);
								data_out(89) <=mem(417)(column_rd_addr);
								data_out(88) <=mem(416)(column_rd_addr);
								data_out(103) <=mem(415)(column_rd_addr);
								data_out(102) <=mem(414)(column_rd_addr);
								data_out(101) <=mem(413)(column_rd_addr);
								data_out(100) <=mem(412)(column_rd_addr);
								data_out(99) <=mem(411)(column_rd_addr);
								data_out(98) <=mem(410)(column_rd_addr);
								data_out(97) <=mem(409)(column_rd_addr);
								data_out(96) <=mem(408)(column_rd_addr);
								data_out(111) <=mem(407)(column_rd_addr);
								data_out(110) <=mem(406)(column_rd_addr);
								data_out(109) <=mem(405)(column_rd_addr);
								data_out(108) <=mem(404)(column_rd_addr);
								data_out(107) <=mem(403)(column_rd_addr);
								data_out(106) <=mem(402)(column_rd_addr);
								data_out(105) <=mem(401)(column_rd_addr);
								data_out(104) <=mem(400)(column_rd_addr);
								data_out(119) <=mem(399)(column_rd_addr);
								data_out(118) <=mem(398)(column_rd_addr);
								data_out(117) <=mem(397)(column_rd_addr);
								data_out(116) <=mem(396)(column_rd_addr);
								data_out(115) <=mem(395)(column_rd_addr);
								data_out(114) <=mem(394)(column_rd_addr);
								data_out(113) <=mem(393)(column_rd_addr);
								data_out(112) <=mem(392)(column_rd_addr);
								data_out(127) <=mem(391)(column_rd_addr);
								data_out(126) <=mem(390)(column_rd_addr);
								data_out(125) <=mem(389)(column_rd_addr);
								data_out(124) <=mem(388)(column_rd_addr);
								data_out(123) <=mem(387)(column_rd_addr);
								data_out(122) <=mem(386)(column_rd_addr);
								data_out(121) <=mem(385)(column_rd_addr);
								data_out(120) <=mem(384)(column_rd_addr);
								data_out(135) <=mem(383)(column_rd_addr);
								data_out(134) <=mem(382)(column_rd_addr);
								data_out(133) <=mem(381)(column_rd_addr);
								data_out(132) <=mem(380)(column_rd_addr);
								data_out(131) <=mem(379)(column_rd_addr);
								data_out(130) <=mem(378)(column_rd_addr);
								data_out(129) <=mem(377)(column_rd_addr);
								data_out(128) <=mem(376)(column_rd_addr);
								data_out(143) <=mem(375)(column_rd_addr);
								data_out(142) <=mem(374)(column_rd_addr);
								data_out(141) <=mem(373)(column_rd_addr);
								data_out(140) <=mem(372)(column_rd_addr);
								data_out(139) <=mem(371)(column_rd_addr);
								data_out(138) <=mem(370)(column_rd_addr);
								data_out(137) <=mem(369)(column_rd_addr);
								data_out(136) <=mem(368)(column_rd_addr);
								data_out(151) <=mem(367)(column_rd_addr);
								data_out(150) <=mem(366)(column_rd_addr);
								data_out(149) <=mem(365)(column_rd_addr);
								data_out(148) <=mem(364)(column_rd_addr);
								data_out(147) <=mem(363)(column_rd_addr);
								data_out(146) <=mem(362)(column_rd_addr);
								data_out(145) <=mem(361)(column_rd_addr);
								data_out(144) <=mem(360)(column_rd_addr);
								data_out(159) <=mem(359)(column_rd_addr);
								data_out(158) <=mem(358)(column_rd_addr);
								data_out(157) <=mem(357)(column_rd_addr);
								data_out(156) <=mem(356)(column_rd_addr);
								data_out(155) <=mem(355)(column_rd_addr);
								data_out(154) <=mem(354)(column_rd_addr);
								data_out(153) <=mem(353)(column_rd_addr);
								data_out(152) <=mem(352)(column_rd_addr);
								data_out(167) <=mem(351)(column_rd_addr);
								data_out(166) <=mem(350)(column_rd_addr);
								data_out(165) <=mem(349)(column_rd_addr);
								data_out(164) <=mem(348)(column_rd_addr);
								data_out(163) <=mem(347)(column_rd_addr);
								data_out(162) <=mem(346)(column_rd_addr);
								data_out(161) <=mem(345)(column_rd_addr);
								data_out(160) <=mem(344)(column_rd_addr);
								data_out(175) <=mem(343)(column_rd_addr);
								data_out(174) <=mem(342)(column_rd_addr);
								data_out(173) <=mem(341)(column_rd_addr);
								data_out(172) <=mem(340)(column_rd_addr);
								data_out(171) <=mem(339)(column_rd_addr);
								data_out(170) <=mem(338)(column_rd_addr);
								data_out(169) <=mem(337)(column_rd_addr);
								data_out(168) <=mem(336)(column_rd_addr);
								data_out(183) <=mem(335)(column_rd_addr);
								data_out(182) <=mem(334)(column_rd_addr);
								data_out(181) <=mem(333)(column_rd_addr);
								data_out(180) <=mem(332)(column_rd_addr);
								data_out(179) <=mem(331)(column_rd_addr);
								data_out(178) <=mem(330)(column_rd_addr);
								data_out(177) <=mem(329)(column_rd_addr);
								data_out(176) <=mem(328)(column_rd_addr);
								data_out(191) <=mem(327)(column_rd_addr);
								data_out(190) <=mem(326)(column_rd_addr);
								data_out(189) <=mem(325)(column_rd_addr);
								data_out(188) <=mem(324)(column_rd_addr);
								data_out(187) <=mem(323)(column_rd_addr);
								data_out(186) <=mem(322)(column_rd_addr);
								data_out(185) <=mem(321)(column_rd_addr);
								data_out(184) <=mem(320)(column_rd_addr);
								data_out(199)<=mem(319)(column_rd_addr);
								data_out(198)<=mem(318)(column_rd_addr);
								data_out(197)<=mem(317)(column_rd_addr);
								data_out(196)<=mem(316)(column_rd_addr);
								data_out(195)<=mem(315)(column_rd_addr);
								data_out(194)<=mem(314)(column_rd_addr);
								data_out(193)<=mem(313)(column_rd_addr);
								data_out(192)<=mem(312)(column_rd_addr);
								data_out(207)<=mem(311)(column_rd_addr);
								data_out(206)<=mem(310)(column_rd_addr);
								data_out(205)<=mem(309)(column_rd_addr);
								data_out(204)<=mem(308)(column_rd_addr);
								data_out(203)<=mem(307)(column_rd_addr);
								data_out(202)<=mem(306)(column_rd_addr);
								data_out(201)<=mem(305)(column_rd_addr);
								data_out(200)<=mem(304)(column_rd_addr);
								data_out(215)<=mem(303)(column_rd_addr);
								data_out(214)<=mem(302)(column_rd_addr);
								data_out(213)<=mem(301)(column_rd_addr);
								data_out(212)<=mem(300)(column_rd_addr);
								data_out(211)<=mem(299)(column_rd_addr);
								data_out(210)<=mem(298)(column_rd_addr);
								data_out(209)<=mem(297)(column_rd_addr);
								data_out(208)<=mem(296)(column_rd_addr);
								data_out(223)<=mem(295)(column_rd_addr);
								data_out(222)<=mem(294)(column_rd_addr);
								data_out(221)<=mem(293)(column_rd_addr);
								data_out(220)<=mem(292)(column_rd_addr);
								data_out(219)<=mem(291)(column_rd_addr);
								data_out(218)<=mem(290)(column_rd_addr);
								data_out(217)<=mem(289)(column_rd_addr);
								data_out(216)<=mem(288)(column_rd_addr);
								data_out(231)<=mem(287)(column_rd_addr);
								data_out(230)<=mem(286)(column_rd_addr);
								data_out(229)<=mem(285)(column_rd_addr);
								data_out(228)<=mem(284)(column_rd_addr);
								data_out(227)<=mem(283)(column_rd_addr);
								data_out(226)<=mem(282)(column_rd_addr);
								data_out(225)<=mem(281)(column_rd_addr);
								data_out(224)<=mem(280)(column_rd_addr);
								data_out(239)<=mem(279)(column_rd_addr);
								data_out(238)<=mem(278)(column_rd_addr);
								data_out(237)<=mem(277)(column_rd_addr);
								data_out(236)<=mem(276)(column_rd_addr);
								data_out(235)<=mem(275)(column_rd_addr);
								data_out(234)<=mem(274)(column_rd_addr);
								data_out(233)<=mem(273)(column_rd_addr);
								data_out(232)<=mem(272)(column_rd_addr);
								data_out(247)<=mem(271)(column_rd_addr);
								data_out(246)<=mem(270)(column_rd_addr);
								data_out(245)<=mem(269)(column_rd_addr);
								data_out(244)<=mem(268)(column_rd_addr);
								data_out(243)<=mem(267)(column_rd_addr);
								data_out(242)<=mem(266)(column_rd_addr);
								data_out(241)<=mem(265)(column_rd_addr);
								data_out(240)<=mem(264)(column_rd_addr);
								data_out(255)<=mem(263)(column_rd_addr);
								data_out(254)<=mem(262)(column_rd_addr);
								data_out(253)<=mem(261)(column_rd_addr);
								data_out(252)<=mem(260)(column_rd_addr);
								data_out(251)<=mem(259)(column_rd_addr);
								data_out(250)<=mem(258)(column_rd_addr);
								data_out(249)<=mem(257)(column_rd_addr);
								data_out(248)<=mem(256)(column_rd_addr);
								data_out(263)<=mem(255)(column_rd_addr);
								data_out(262)<=mem(254)(column_rd_addr);
								data_out(261)<=mem(253)(column_rd_addr);
								data_out(260)<=mem(252)(column_rd_addr);
								data_out(259)<=mem(251)(column_rd_addr);
								data_out(258)<=mem(250)(column_rd_addr);
								data_out(257)<=mem(249)(column_rd_addr);
								data_out(256)<=mem(248)(column_rd_addr);
								data_out(271)<=mem(247)(column_rd_addr);
								data_out(270)<=mem(246)(column_rd_addr);
								data_out(269)<=mem(245)(column_rd_addr);
								data_out(268)<=mem(244)(column_rd_addr);
								data_out(267)<=mem(243)(column_rd_addr);
								data_out(266)<=mem(242)(column_rd_addr);
								data_out(265)<=mem(241)(column_rd_addr);
								data_out(264)<=mem(240)(column_rd_addr);
								data_out(279)<=mem(239)(column_rd_addr);
								data_out(278)<=mem(238)(column_rd_addr);
								data_out(277)<=mem(237)(column_rd_addr);
								data_out(276)<=mem(236)(column_rd_addr);
								data_out(275)<=mem(235)(column_rd_addr);
								data_out(274)<=mem(234)(column_rd_addr);
								data_out(273)<=mem(233)(column_rd_addr);
								data_out(272)<=mem(232)(column_rd_addr);
								data_out(287)<=mem(231)(column_rd_addr);
								data_out(286)<=mem(230)(column_rd_addr);
								data_out(285)<=mem(229)(column_rd_addr);
								data_out(284)<=mem(228)(column_rd_addr);
								data_out(283)<=mem(227)(column_rd_addr);
								data_out(282)<=mem(226)(column_rd_addr);
								data_out(281)<=mem(225)(column_rd_addr);
								data_out(280)<=mem(224)(column_rd_addr);
								data_out(295)<=mem(223)(column_rd_addr);
								data_out(294)<=mem(222)(column_rd_addr);
								data_out(293)<=mem(221)(column_rd_addr);
								data_out(292)<=mem(220)(column_rd_addr);
								data_out(291)<=mem(219)(column_rd_addr);
								data_out(290)<=mem(218)(column_rd_addr);
								data_out(289)<=mem(217)(column_rd_addr);
								data_out(288)<=mem(216)(column_rd_addr);
								data_out(303)<=mem(215)(column_rd_addr);
								data_out(302)<=mem(214)(column_rd_addr);
								data_out(301)<=mem(213)(column_rd_addr);
								data_out(300)<=mem(212)(column_rd_addr);
								data_out(299)<=mem(211)(column_rd_addr);
								data_out(298)<=mem(210)(column_rd_addr);
								data_out(297)<=mem(209)(column_rd_addr);
								data_out(296)<=mem(208)(column_rd_addr);
								data_out(311)<=mem(207)(column_rd_addr);
								data_out(310)<=mem(206)(column_rd_addr);
								data_out(309)<=mem(205)(column_rd_addr);
								data_out(308)<=mem(204)(column_rd_addr);
								data_out(307)<=mem(203)(column_rd_addr);
								data_out(306)<=mem(202)(column_rd_addr);
								data_out(305)<=mem(201)(column_rd_addr);
								data_out(304)<=mem(200)(column_rd_addr);
								data_out(319)<=mem(199)(column_rd_addr);
								data_out(318)<=mem(198)(column_rd_addr);
								data_out(317)<=mem(197)(column_rd_addr);
								data_out(316)<=mem(196)(column_rd_addr);
								data_out(315)<=mem(195)(column_rd_addr);
								data_out(314)<=mem(194)(column_rd_addr);
								data_out(313)<=mem(193)(column_rd_addr);
								data_out(312)<=mem(192)(column_rd_addr);
								data_out(327)<=mem(191)(column_rd_addr);
								data_out(326)<=mem(190)(column_rd_addr);
								data_out(325)<=mem(189)(column_rd_addr);
								data_out(324)<=mem(188)(column_rd_addr);
								data_out(323)<=mem(187)(column_rd_addr);
								data_out(322)<=mem(186)(column_rd_addr);
								data_out(321)<=mem(185)(column_rd_addr);
								data_out(320)<=mem(184)(column_rd_addr);
								data_out(335)<=mem(183)(column_rd_addr);
								data_out(334)<=mem(182)(column_rd_addr);
								data_out(333)<=mem(181)(column_rd_addr);
								data_out(332)<=mem(180)(column_rd_addr);
								data_out(331)<=mem(179)(column_rd_addr);
								data_out(330)<=mem(178)(column_rd_addr);
								data_out(329)<=mem(177)(column_rd_addr);
								data_out(328)<=mem(176)(column_rd_addr);
								data_out(343)<=mem(175)(column_rd_addr);
								data_out(342)<=mem(174)(column_rd_addr);
								data_out(341)<=mem(173)(column_rd_addr);
								data_out(340)<=mem(172)(column_rd_addr);
								data_out(339)<=mem(171)(column_rd_addr);
								data_out(338)<=mem(170)(column_rd_addr);
								data_out(337)<=mem(169)(column_rd_addr);
								data_out(336)<=mem(168)(column_rd_addr);
								data_out(351)<=mem(167)(column_rd_addr);
								data_out(350)<=mem(166)(column_rd_addr);
								data_out(349)<=mem(165)(column_rd_addr);
								data_out(348)<=mem(164)(column_rd_addr);
								data_out(347)<=mem(163)(column_rd_addr);
								data_out(346)<=mem(162)(column_rd_addr);
								data_out(345)<=mem(161)(column_rd_addr);
								data_out(344)<=mem(160)(column_rd_addr);
								data_out(359)<=mem(159)(column_rd_addr);
								data_out(358)<=mem(158)(column_rd_addr);
								data_out(357)<=mem(157)(column_rd_addr);
								data_out(356)<=mem(156)(column_rd_addr);
								data_out(355)<=mem(155)(column_rd_addr);
								data_out(354)<=mem(154)(column_rd_addr);
								data_out(353)<=mem(153)(column_rd_addr);
								data_out(352)<=mem(152)(column_rd_addr);
								data_out(367)<=mem(151)(column_rd_addr);
								data_out(366)<=mem(150)(column_rd_addr);
								data_out(365)<=mem(149)(column_rd_addr);
								data_out(364)<=mem(148)(column_rd_addr);
								data_out(363)<=mem(147)(column_rd_addr);
								data_out(362)<=mem(146)(column_rd_addr);
								data_out(361)<=mem(145)(column_rd_addr);
								data_out(360)<=mem(144)(column_rd_addr);
								data_out(375)<=mem(143)(column_rd_addr);
								data_out(374)<=mem(142)(column_rd_addr);
								data_out(373)<=mem(141)(column_rd_addr);
								data_out(372)<=mem(140)(column_rd_addr);
								data_out(371)<=mem(139)(column_rd_addr);
								data_out(370)<=mem(138)(column_rd_addr);
								data_out(369)<=mem(137)(column_rd_addr);
								data_out(368)<=mem(136)(column_rd_addr);
								data_out(383)<=mem(135)(column_rd_addr);
								data_out(382)<=mem(134)(column_rd_addr);
								data_out(381)<=mem(133)(column_rd_addr);
								data_out(380)<=mem(132)(column_rd_addr);
								data_out(379)<=mem(131)(column_rd_addr);
								data_out(378)<=mem(130)(column_rd_addr);
								data_out(377)<=mem(129)(column_rd_addr);
								data_out(376)<=mem(128)(column_rd_addr);
								data_out(391)<=mem(127)(column_rd_addr);
								data_out(390)<=mem(126)(column_rd_addr);
								data_out(389)<=mem(125)(column_rd_addr);
								data_out(388)<=mem(124)(column_rd_addr);
								data_out(387)<=mem(123)(column_rd_addr);
								data_out(386)<=mem(122)(column_rd_addr);
								data_out(385)<=mem(121)(column_rd_addr);
								data_out(384)<=mem(120)(column_rd_addr);
								data_out(399)<=mem(119)(column_rd_addr);
								data_out(398)<=mem(118)(column_rd_addr);
								data_out(397)<=mem(117)(column_rd_addr);
								data_out(396)<=mem(116)(column_rd_addr);
								data_out(395)<=mem(115)(column_rd_addr);
								data_out(394)<=mem(114)(column_rd_addr);
								data_out(393)<=mem(113)(column_rd_addr);
								data_out(392)<=mem(112)(column_rd_addr);
								data_out(407)<=mem(111)(column_rd_addr);
								data_out(406)<=mem(110)(column_rd_addr);
								data_out(405)<=mem(109)(column_rd_addr);
								data_out(404)<=mem(108)(column_rd_addr);
								data_out(403)<=mem(107)(column_rd_addr);
								data_out(402)<=mem(106)(column_rd_addr);
								data_out(401)<=mem(105)(column_rd_addr);
								data_out(400)<=mem(104)(column_rd_addr);
								data_out(415)<=mem(103)(column_rd_addr);
								data_out(414)<=mem(102)(column_rd_addr);
								data_out(413)<=mem(101)(column_rd_addr);
								data_out(412)<=mem(100)(column_rd_addr);
								data_out(411)<=mem(99)(column_rd_addr);
								data_out(410)<=mem(98)(column_rd_addr);
								data_out(409)<=mem(97)(column_rd_addr);
								data_out(408)<=mem(96)(column_rd_addr);
								data_out(423)<=mem(95)(column_rd_addr);
								data_out(422)<=mem(94)(column_rd_addr);
								data_out(421)<=mem(93)(column_rd_addr);
								data_out(420)<=mem(92)(column_rd_addr);
								data_out(419)<=mem(91)(column_rd_addr);
								data_out(418)<=mem(90)(column_rd_addr);
								data_out(417)<=mem(89)(column_rd_addr);
								data_out(416)<=mem(88)(column_rd_addr);
								data_out(431)<=mem(87)(column_rd_addr);
								data_out(430)<=mem(86)(column_rd_addr);
								data_out(429)<=mem(85)(column_rd_addr);
								data_out(428)<=mem(84)(column_rd_addr);
								data_out(427)<=mem(83)(column_rd_addr);
								data_out(426)<=mem(82)(column_rd_addr);
								data_out(425)<=mem(81)(column_rd_addr);
								data_out(424)<=mem(80)(column_rd_addr);
								data_out(439)<=mem(79)(column_rd_addr);
								data_out(438)<=mem(78)(column_rd_addr);
								data_out(437)<=mem(77)(column_rd_addr);
								data_out(436)<=mem(76)(column_rd_addr);
								data_out(435)<=mem(75)(column_rd_addr);
								data_out(434)<=mem(74)(column_rd_addr);
								data_out(433)<=mem(73)(column_rd_addr);
								data_out(432)<=mem(72)(column_rd_addr);
								data_out(447)<=mem(71)(column_rd_addr);
								data_out(446)<=mem(70)(column_rd_addr);
								data_out(445)<=mem(69)(column_rd_addr);
								data_out(444)<=mem(68)(column_rd_addr);
								data_out(443)<=mem(67)(column_rd_addr);
								data_out(442)<=mem(66)(column_rd_addr);
								data_out(441)<=mem(65)(column_rd_addr);
								data_out(440)<=mem(64)(column_rd_addr);
								data_out(455)<=mem(63)(column_rd_addr);
								data_out(454)<=mem(62)(column_rd_addr);
								data_out(453)<=mem(61)(column_rd_addr);
								data_out(452)<=mem(60)(column_rd_addr);
								data_out(451)<=mem(59)(column_rd_addr);
								data_out(450)<=mem(58)(column_rd_addr);
								data_out(449)<=mem(57)(column_rd_addr);
								data_out(448)<=mem(56)(column_rd_addr);
								data_out(463)<=mem(55)(column_rd_addr);
								data_out(462)<=mem(54)(column_rd_addr);
								data_out(461)<=mem(53)(column_rd_addr);
								data_out(460)<=mem(52)(column_rd_addr);
								data_out(459)<=mem(51)(column_rd_addr);
								data_out(458)<=mem(50)(column_rd_addr);
								data_out(457)<=mem(49)(column_rd_addr);
								data_out(456)<=mem(48)(column_rd_addr);
								data_out(471)<=mem(47)(column_rd_addr);
								data_out(470)<=mem(46)(column_rd_addr);
								data_out(469)<=mem(45)(column_rd_addr);
								data_out(468)<=mem(44)(column_rd_addr);
								data_out(467)<=mem(43)(column_rd_addr);
								data_out(466)<=mem(42)(column_rd_addr);
								data_out(465)<=mem(41)(column_rd_addr);
								data_out(464)<=mem(40)(column_rd_addr);
								data_out(479)<=mem(39)(column_rd_addr);
								data_out(478)<=mem(38)(column_rd_addr);
								data_out(477)<=mem(37)(column_rd_addr);
								data_out(476)<=mem(36)(column_rd_addr);
								data_out(475)<=mem(35)(column_rd_addr);
								data_out(474)<=mem(34)(column_rd_addr);
								data_out(473)<=mem(33)(column_rd_addr);
								data_out(472)<=mem(32)(column_rd_addr);
								data_out(487)<=mem(31)(column_rd_addr);
								data_out(486)<=mem(30)(column_rd_addr);
								data_out(485)<=mem(29)(column_rd_addr);
								data_out(484)<=mem(28)(column_rd_addr);
								data_out(483)<=mem(27)(column_rd_addr);
								data_out(482)<=mem(26)(column_rd_addr);
								data_out(481)<=mem(25)(column_rd_addr);
								data_out(480)<=mem(24)(column_rd_addr);
								data_out(495)<=mem(23)(column_rd_addr);
								data_out(494)<=mem(22)(column_rd_addr);
								data_out(493)<=mem(21)(column_rd_addr);
								data_out(492)<=mem(20)(column_rd_addr);
								data_out(491)<=mem(19)(column_rd_addr);
								data_out(490)<=mem(18)(column_rd_addr);
								data_out(489)<=mem(17)(column_rd_addr);
								data_out(488)<=mem(16)(column_rd_addr);
								data_out(503)<=mem(15)(column_rd_addr);
								data_out(502)<=mem(14)(column_rd_addr);
								data_out(501)<=mem(13)(column_rd_addr);
								data_out(500)<=mem(12)(column_rd_addr);
								data_out(499)<=mem(11)(column_rd_addr);
								data_out(498)<=mem(10)(column_rd_addr);
								data_out(497)<=mem(9)(column_rd_addr);
								data_out(496)<=mem(8)(column_rd_addr);
								data_out(511)<=mem(7)(column_rd_addr);
								data_out(510)<=mem(6)(column_rd_addr);
								data_out(509)<=mem(5)(column_rd_addr);
								data_out(508)<=mem(4)(column_rd_addr);
								data_out(507)<=mem(3)(column_rd_addr);
								data_out(506)<=mem(2)(column_rd_addr);
								data_out(505)<=mem(1)(column_rd_addr);
								data_out(504)<=mem(0)(column_rd_addr);

			END IF;	
	END PROCESS;
END behavioral;